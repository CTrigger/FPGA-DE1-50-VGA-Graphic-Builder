ENTITY Projeto_Base IS
	PORT
	(
		-- INDICANDO QUE SERA USADO O CLOCK DE 27 MHZ
		CLOCK_27 : IN bit_vector (0 to 1);
		CLOCK_50 : IN bit;
		
		-- PINOS DE SAIDA DO SINCRONISMO
		VGA_VS, VGA_HS : BUFFER BIT;
		
		-- Controles de cor
		VGA_R: out integer range 15 downto 0 := 0;
		VGA_G: out integer range 15 downto 0 := 0;
		VGA_B: out integer range 15 downto 0 := 0;
		-- VGA_R: BUFFER bit_vector (0 to 3);
		-- VGA_G: BUFFER bit_vector (0 to 3);
		-- VGA_B: BUFFER bit_vector (0 to 3);
		
		-- leds confirmacao visual
		LEDG: BUFFER bit_vector (0 to 7);
		
		-- botoes de movimento
		KEY: IN bit_vector (0 to 3)
		
	);
END Projeto_Base;
 
ARCHITECTURE Kim OF Projeto_Base IS

	-- controle de clock do video (compensar 27 MHz)
	SIGNAL countHS: integer RANGE 0 TO 809;
	SIGNAL countVS: integer RANGE 0 TO 525;

	-- controle de sinal
	SIGNAL enableHS: bit;
	SIGNAL enableVS: bit;
	
	-- Controle do display
	SIGNAL drawHS: integer RANGE 0 TO 640 := 0;
	SIGNAL drawVS: integer RANGE 0 TO 480 := 0;
	
	SIGNAL showColor: bit;
	SIGNAL hideColor: bit;
	SIGNAL showDisplay: boolean;
	
	-- Controle do desenho
	SIGNAL startController: bit;
	SIGNAL xInit, xEnd: integer RANGE 0 TO 640;
	SIGNAL yInit, yEnd: integer RANGE 0 TO 480;
	SIGNAL quadrado: boolean;
	
	-- Controle de Direcao
	CONSTANT cima: integer := 0;
	CONSTANT baixo: integer := 1;
	CONSTANT esquerda: integer := 2;
	CONSTANT direita: integer := 3;
	CONSTANT tempo: integer := 700000;
	SIGNAL moveDelay: integer RANGE 0 TO tempo;
	
	
	-- ================================
	--            Desenhos
	-- ================================

	--Pacman
	SIGNAL pacmanFrame: integer RANGE 0 TO 3;
	TYPE cor IS
		RECORD
			r: integer RANGE 15 DOWNTO 0;
			g: integer RANGE 15 DOWNTO 0;
			b: integer RANGE 15 DOWNTO 0;
		END RECORD;
	TYPE matriz IS ARRAY(0 TO 9, 0 TO 9) OF cor;
	TYPE frames IS ARRAY(0 TO 3) OF matriz;
	CONSTANT pacman: frames := (
		 0 => (
			0 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)), 
			1 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			2 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			3 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			4 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			5 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			6 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			7 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			8 => (0 => (0,0,15), 1 => (15,15,0), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (15,15,0), 9 => (0,0,15)), 
			9 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)) 
		 ),
		 
		 1 => (
			0 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)), 
			1 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			2 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			3 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			4 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			5 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (0,0,15), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			6 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			7 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			8 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (15,15,0), 9 => (0,0,15)), 
			9 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)) 
		 ),
		 
		 2 => (
			0 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)), 
			1 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			2 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			3 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			4 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			5 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			6 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (0,0,15), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			7 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			8 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			9 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (0,0,15), 4 => (0,0,15), 5 => (0,0,15), 6 => (0,0,15), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)) 

		 ),
		 
		 3 => (
			0 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)), 
			1 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			2 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			3 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			4 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			5 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			6 => (0 => (15,15,0), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (15,15,0)), 
			7 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			8 => (0 => (0,0,15), 1 => (15,15,0), 2 => (15,15,0), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (15,15,0), 8 => (15,15,0), 9 => (0,0,15)), 
			9 => (0 => (0,0,15), 1 => (0,0,15), 2 => (0,0,15), 3 => (15,15,0), 4 => (15,15,0), 5 => (15,15,0), 6 => (15,15,0), 7 => (0,0,15), 8 => (0,0,15), 9 => (0,0,15)) 
		)
	);
	
	--SONIC BACKGROUND
	SIGNAL sonicBG: integer RANGE 0 TO 0;
	TYPE sonicMatriz IS ARRAY(0 TO 111, 0 TO 159) OF cor;
	TYPE sonicFrames IS ARRAY(0 TO 0) OF sonicMatriz;
	CONSTANT sonic: sonicFrames := (
		0 => (
			0 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			1 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			2 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			3 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			4 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			5 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			6 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			7 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			8 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			9 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			10 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			11 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			12 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			13 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			14 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			15 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			16 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,1,14), 18 => (0,1,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,1,14), 73 => (0,1,14), 74 => (0,1,14), 75 => (0,1,14), 76 => (0,1,14), 77 => (0,1,14), 78 => (0,1,14), 79 => (0,1,14), 80 => (0,1,14), 81 => (0,1,14), 82 => (0,1,14), 83 => (0,1,14), 84 => (0,1,14), 85 => (0,1,14), 86 => (0,1,14), 87 => (0,1,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,15), 98 => (0,0,12), 99 => (0,0,12), 100 => (0,0,12), 101 => (0,0,12), 102 => (0,0,12), 103 => (0,1,13), 104 => (0,1,14), 105 => (0,1,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,1,14), 142 => (0,1,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			17 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (1,1,8), 17 => (4,4,8), 18 => (4,5,15), 19 => (0,0,8), 20 => (0,1,14), 21 => (0,1,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,1,14), 69 => (0,1,14), 70 => (0,1,14), 71 => (0,0,13), 72 => (5,6,14), 73 => (8,9,14), 74 => (10,9,13), 75 => (10,10,14), 76 => (10,10,14), 77 => (10,10,14), 78 => (10,10,14), 79 => (10,10,14), 80 => (10,10,14), 81 => (10,10,14), 82 => (10,10,14), 83 => (10,10,14), 84 => (10,10,14), 85 => (10,9,13), 86 => (8,9,14), 87 => (5,6,14), 88 => (0,0,13), 89 => (0,1,14), 90 => (0,1,14), 91 => (0,1,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,0,12), 95 => (1,1,12), 96 => (1,1,13), 97 => (0,0,2), 98 => (4,3,15), 99 => (3,3,14), 100 => (3,3,14), 101 => (3,3,14), 102 => (3,3,14), 103 => (3,3,14), 104 => (3,3,14), 105 => (2,2,14), 106 => (0,1,14), 107 => (0,1,14), 108 => (0,1,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,1,14), 139 => (0,1,14), 140 => (0,0,8), 141 => (4,5,15), 142 => (4,4,8), 143 => (1,1,8), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			18 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,0,4), 17 => (6,5,14), 18 => (12,12,14), 19 => (14,13,14), 20 => (6,5,13), 21 => (3,3,9), 22 => (0,0,8), 23 => (0,1,14), 24 => (0,1,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,1,14), 67 => (0,1,14), 68 => (0,1,13), 69 => (8,8,13), 70 => (11,11,14), 71 => (10,10,14), 72 => (7,7,14), 73 => (4,4,14), 74 => (5,5,14), 75 => (7,7,15), 76 => (7,7,15), 77 => (7,7,15), 78 => (7,7,15), 79 => (7,7,15), 80 => (7,7,15), 81 => (7,7,15), 82 => (7,7,15), 83 => (7,7,15), 84 => (7,7,15), 85 => (5,5,14), 86 => (4,4,14), 87 => (7,7,14), 88 => (10,10,14), 89 => (11,11,14), 90 => (8,9,13), 91 => (1,2,13), 92 => (0,0,12), 93 => (2,1,12), 94 => (5,5,14), 95 => (1,1,14), 96 => (5,6,14), 97 => (6,6,15), 98 => (0,0,3), 99 => (2,2,15), 100 => (1,1,14), 101 => (1,1,14), 102 => (1,1,14), 103 => (1,1,14), 104 => (1,1,14), 105 => (2,2,14), 106 => (3,3,14), 107 => (3,3,14), 108 => (2,2,14), 109 => (0,0,12), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,1,14), 136 => (0,1,14), 137 => (0,0,8), 138 => (3,3,9), 139 => (6,5,13), 140 => (14,13,14), 141 => (12,12,14), 142 => (6,5,14), 143 => (0,0,4), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			19 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,0,4), 17 => (2,2,14), 18 => (10,10,14), 19 => (15,15,14), 20 => (15,15,14), 21 => (14,13,14), 22 => (13,13,14), 23 => (6,5,13), 24 => (3,3,9), 25 => (0,0,8), 26 => (0,1,14), 27 => (0,1,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,1,14), 65 => (0,0,13), 66 => (5,5,13), 67 => (11,11,14), 68 => (10,10,14), 69 => (4,4,14), 70 => (5,5,14), 71 => (7,7,15), 72 => (4,4,14), 73 => (2,3,14), 74 => (3,4,15), 75 => (4,1,4), 76 => (4,2,5), 77 => (4,2,5), 78 => (4,2,5), 79 => (4,2,5), 80 => (4,2,5), 81 => (4,2,5), 82 => (4,2,5), 83 => (4,2,5), 84 => (4,1,4), 85 => (3,4,15), 86 => (2,3,14), 87 => (4,4,14), 88 => (8,8,14), 89 => (3,3,13), 90 => (0,0,12), 91 => (3,3,13), 92 => (4,4,14), 93 => (2,2,14), 94 => (1,1,14), 95 => (5,6,14), 96 => (3,2,11), 97 => (4,2,7), 98 => (0,1,11), 99 => (1,1,10), 100 => (2,2,14), 101 => (2,2,14), 102 => (2,2,14), 103 => (2,2,14), 104 => (2,2,14), 105 => (1,1,14), 106 => (1,1,14), 107 => (1,1,14), 108 => (3,3,14), 109 => (3,3,14), 110 => (2,2,12), 111 => (0,0,12), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,1,14), 133 => (0,1,14), 134 => (0,0,8), 135 => (3,3,9), 136 => (6,5,13), 137 => (13,13,14), 138 => (14,13,14), 139 => (15,15,14), 140 => (15,15,14), 141 => (10,10,14), 142 => (2,2,14), 143 => (0,0,4), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			20 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,15), 17 => (0,0,3), 18 => (8,8,15), 19 => (12,12,14), 20 => (14,14,14), 21 => (14,14,14), 22 => (14,14,14), 23 => (15,15,14), 24 => (14,13,14), 25 => (13,13,14), 26 => (6,5,13), 27 => (3,3,9), 28 => (0,0,8), 29 => (0,1,14), 30 => (0,1,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,1,14), 63 => (0,0,13), 64 => (5,5,13), 65 => (12,11,14), 66 => (7,7,14), 67 => (4,4,14), 68 => (7,7,14), 69 => (4,4,14), 70 => (3,4,15), 71 => (3,1,5), 72 => (9,6,2), 73 => (11,6,0), 74 => (10,6,0), 75 => (10,5,0), 76 => (10,5,0), 77 => (10,5,0), 78 => (10,5,0), 79 => (10,5,0), 80 => (10,5,0), 81 => (10,5,0), 82 => (10,5,0), 83 => (10,5,0), 84 => (10,5,0), 85 => (10,6,0), 86 => (11,6,0), 87 => (7,4,4), 88 => (0,0,12), 89 => (4,4,13), 90 => (6,6,14), 91 => (2,2,14), 92 => (1,1,14), 93 => (1,1,14), 94 => (5,5,14), 95 => (2,2,12), 96 => (9,5,0), 97 => (11,6,2), 98 => (3,3,12), 99 => (0,0,3), 100 => (2,2,15), 101 => (2,2,14), 102 => (2,2,14), 103 => (2,2,14), 104 => (2,2,14), 105 => (2,2,14), 106 => (2,2,14), 107 => (2,2,14), 108 => (1,1,14), 109 => (1,1,14), 110 => (2,2,14), 111 => (2,2,14), 112 => (1,0,12), 113 => (0,0,13), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,1,14), 130 => (0,1,14), 131 => (0,0,8), 132 => (3,3,9), 133 => (6,5,13), 134 => (13,13,14), 135 => (14,13,14), 136 => (15,15,14), 137 => (14,14,14), 138 => (14,14,14), 139 => (14,14,14), 140 => (12,12,14), 141 => (8,8,15), 142 => (0,0,3), 143 => (0,2,15), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			21 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,0,4), 18 => (2,2,14), 19 => (10,10,14), 20 => (14,14,14), 21 => (14,14,14), 22 => (14,14,14), 23 => (14,14,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (15,15,14), 27 => (14,13,14), 28 => (13,13,14), 29 => (6,5,13), 30 => (3,3,9), 31 => (0,0,8), 32 => (0,1,14), 33 => (0,1,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,0,13), 62 => (5,6,13), 63 => (10,10,14), 64 => (7,7,14), 65 => (4,4,14), 66 => (7,7,14), 67 => (4,4,15), 68 => (3,3,11), 69 => (9,6,2), 70 => (10,5,0), 71 => (10,5,0), 72 => (11,7,0), 73 => (5,6,15), 74 => (10,7,3), 75 => (15,13,0), 76 => (14,12,0), 77 => (14,12,0), 78 => (14,12,0), 79 => (14,12,0), 80 => (14,12,0), 81 => (14,12,0), 82 => (14,12,0), 83 => (14,12,0), 84 => (15,13,0), 85 => (11,7,2), 86 => (4,4,11), 87 => (2,2,14), 88 => (6,6,14), 89 => (4,4,14), 90 => (1,1,14), 91 => (1,1,14), 92 => (1,1,14), 93 => (4,4,14), 94 => (4,4,12), 95 => (9,4,0), 96 => (12,8,6), 97 => (12,8,5), 98 => (5,3,8), 99 => (0,0,5), 100 => (0,0,13), 101 => (2,2,14), 102 => (2,2,14), 103 => (2,2,14), 104 => (2,2,14), 105 => (2,2,14), 106 => (2,2,14), 107 => (2,2,14), 108 => (2,2,14), 109 => (2,2,14), 110 => (1,1,13), 111 => (0,0,13), 112 => (1,1,14), 113 => (0,0,7), 114 => (0,1,9), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,1,14), 127 => (0,1,14), 128 => (0,0,8), 129 => (3,3,9), 130 => (6,5,13), 131 => (13,13,14), 132 => (14,13,14), 133 => (15,15,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (14,14,14), 137 => (14,14,14), 138 => (14,14,14), 139 => (14,14,14), 140 => (10,10,14), 141 => (2,2,14), 142 => (0,0,4), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			22 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,15), 18 => (0,0,3), 19 => (5,5,14), 20 => (12,12,14), 21 => (14,14,14), 22 => (14,14,14), 23 => (14,14,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (15,15,14), 30 => (14,13,14), 31 => (13,13,14), 32 => (6,5,13), 33 => (3,3,9), 34 => (0,0,8), 35 => (0,1,14), 36 => (0,1,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,1,14), 60 => (0,1,13), 61 => (9,9,13), 62 => (5,5,14), 63 => (4,4,14), 64 => (7,7,14), 65 => (4,4,15), 66 => (3,3,11), 67 => (9,6,2), 68 => (10,5,0), 69 => (11,6,0), 70 => (12,8,0), 71 => (13,10,0), 72 => (12,7,0), 73 => (13,6,0), 74 => (8,3,0), 75 => (7,8,5), 76 => (14,14,0), 77 => (14,14,0), 78 => (14,14,0), 79 => (14,14,0), 80 => (14,14,0), 81 => (14,14,0), 82 => (14,14,0), 83 => (14,14,0), 84 => (9,9,2), 85 => (2,3,9), 86 => (2,3,14), 87 => (6,6,14), 88 => (1,1,14), 89 => (1,1,14), 90 => (2,2,14), 91 => (1,1,14), 92 => (2,2,14), 93 => (5,4,11), 94 => (9,4,0), 95 => (12,8,6), 96 => (13,9,7), 97 => (14,10,8), 98 => (11,6,2), 99 => (1,2,11), 100 => (0,0,8), 101 => (0,0,12), 102 => (1,1,13), 103 => (2,2,14), 104 => (2,2,14), 105 => (1,1,13), 106 => (1,1,13), 107 => (0,0,11), 108 => (0,0,11), 109 => (0,0,11), 110 => (0,0,12), 111 => (0,0,8), 112 => (0,0,3), 113 => (0,1,10), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,1,14), 124 => (0,1,14), 125 => (0,0,8), 126 => (3,3,9), 127 => (6,5,13), 128 => (13,13,14), 129 => (14,13,14), 130 => (15,15,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (14,14,14), 137 => (14,14,14), 138 => (14,14,14), 139 => (12,12,14), 140 => (5,5,14), 141 => (0,0,3), 142 => (0,2,15), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			23 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,1,10), 19 => (0,0,8), 20 => (10,10,15), 21 => (13,13,14), 22 => (14,14,14), 23 => (14,14,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (15,15,14), 33 => (14,13,14), 34 => (13,13,14), 35 => (6,5,13), 36 => (3,3,9), 37 => (0,0,8), 38 => (0,1,14), 39 => (0,1,14), 40 => (0,1,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,1,14), 59 => (0,0,12), 60 => (9,9,14), 61 => (3,3,14), 62 => (7,7,14), 63 => (5,5,15), 64 => (3,2,11), 65 => (9,6,2), 66 => (10,5,0), 67 => (12,7,0), 68 => (13,10,0), 69 => (13,11,0), 70 => (12,8,0), 71 => (11,4,0), 72 => (7,2,1), 73 => (4,0,2), 74 => (10,3,0), 75 => (10,11,0), 76 => (14,15,0), 77 => (14,14,0), 78 => (14,14,0), 79 => (14,14,0), 80 => (14,15,0), 81 => (15,15,0), 82 => (15,15,0), 83 => (15,15,0), 84 => (2,2,10), 85 => (4,4,15), 86 => (4,4,14), 87 => (2,2,14), 88 => (1,1,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (1,1,14), 92 => (2,2,14), 93 => (3,2,10), 94 => (7,5,10), 95 => (11,8,8), 96 => (15,11,7), 97 => (14,10,8), 98 => (11,7,3), 99 => (2,2,15), 100 => (0,0,3), 101 => (0,0,12), 102 => (0,0,11), 103 => (0,0,11), 104 => (0,0,11), 105 => (0,0,11), 106 => (0,0,11), 107 => (0,0,12), 108 => (0,0,12), 109 => (0,0,13), 110 => (0,0,2), 111 => (0,1,10), 112 => (0,2,15), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,1,14), 120 => (0,1,14), 121 => (0,1,14), 122 => (0,0,8), 123 => (3,3,9), 124 => (6,5,13), 125 => (13,13,14), 126 => (14,13,14), 127 => (15,15,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (14,14,14), 137 => (14,14,14), 138 => (13,13,14), 139 => (10,10,15), 140 => (0,0,8), 141 => (0,1,10), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			24 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,1,9), 20 => (0,0,8), 21 => (9,9,14), 22 => (13,13,14), 23 => (14,14,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (15,15,14), 36 => (14,13,14), 37 => (13,13,14), 38 => (11,10,14), 39 => (4,3,8), 40 => (3,4,15), 41 => (0,0,8), 42 => (0,1,14), 43 => (0,1,14), 44 => (0,1,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,1,14), 52 => (0,1,15), 53 => (0,1,15), 54 => (0,2,15), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,0,13), 58 => (6,6,13), 59 => (8,8,14), 60 => (4,4,14), 61 => (8,8,14), 62 => (2,3,15), 63 => (7,3,1), 64 => (10,5,0), 65 => (10,5,0), 66 => (14,12,0), 67 => (14,15,0), 68 => (12,12,0), 69 => (13,8,3), 70 => (13,5,0), 71 => (4,4,9), 72 => (6,9,14), 73 => (5,2,4), 74 => (10,2,0), 75 => (10,12,10), 76 => (12,8,0), 77 => (12,8,0), 78 => (11,7,0), 79 => (11,8,0), 80 => (9,5,0), 81 => (0,0,0), 82 => (0,0,0), 83 => (0,0,1), 84 => (4,4,15), 85 => (4,4,14), 86 => (1,1,14), 87 => (1,1,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (2,2,14), 92 => (1,1,14), 93 => (1,1,14), 94 => (1,1,14), 95 => (0,1,14), 96 => (3,3,13), 97 => (12,9,9), 98 => (12,7,3), 99 => (2,2,15), 100 => (1,1,5), 101 => (0,0,12), 102 => (0,0,12), 103 => (0,0,12), 104 => (0,0,12), 105 => (0,0,12), 106 => (0,0,12), 107 => (0,0,13), 108 => (0,0,4), 109 => (0,0,0), 110 => (0,2,15), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,1,14), 116 => (0,1,14), 117 => (0,1,14), 118 => (0,0,8), 119 => (3,4,15), 120 => (4,3,8), 121 => (11,10,14), 122 => (13,13,14), 123 => (14,13,14), 124 => (15,15,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (14,14,14), 137 => (13,13,14), 138 => (9,9,14), 139 => (0,0,8), 140 => (0,1,9), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			25 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,15), 20 => (0,0,3), 21 => (5,5,15), 22 => (11,11,14), 23 => (14,14,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (15,15,14), 40 => (14,13,14), 41 => (13,13,14), 42 => (11,10,14), 43 => (4,3,8), 44 => (3,4,15), 45 => (0,0,8), 46 => (0,1,14), 47 => (0,1,14), 48 => (0,1,14), 49 => (0,2,14), 50 => (0,1,14), 51 => (5,2,5), 52 => (12,8,5), 53 => (9,3,0), 54 => (8,1,0), 55 => (1,0,7), 56 => (1,0,6), 57 => (5,4,10), 58 => (5,6,15), 59 => (5,6,15), 60 => (5,6,15), 61 => (3,2,11), 62 => (11,6,0), 63 => (11,7,0), 64 => (13,11,0), 65 => (14,14,0), 66 => (14,15,0), 67 => (12,11,0), 68 => (13,9,6), 69 => (12,6,0), 70 => (7,8,13), 71 => (10,12,15), 72 => (8,11,15), 73 => (6,3,6), 74 => (12,6,0), 75 => (12,6,0), 76 => (9,2,0), 77 => (9,6,0), 78 => (14,15,0), 79 => (15,15,0), 80 => (0,0,15), 81 => (0,0,14), 82 => (0,0,0), 83 => (4,4,15), 84 => (4,4,14), 85 => (1,1,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (2,2,14), 92 => (2,2,14), 93 => (2,2,14), 94 => (2,2,14), 95 => (2,2,14), 96 => (1,1,14), 97 => (0,0,15), 98 => (9,5,3), 99 => (2,3,15), 100 => (0,0,4), 101 => (0,0,12), 102 => (0,0,12), 103 => (0,0,12), 104 => (0,0,12), 105 => (0,0,13), 106 => (0,0,10), 107 => (0,0,0), 108 => (0,1,11), 109 => (0,2,15), 110 => (0,2,14), 111 => (0,1,14), 112 => (0,1,14), 113 => (0,1,14), 114 => (0,0,8), 115 => (3,4,15), 116 => (4,3,8), 117 => (11,10,14), 118 => (13,13,14), 119 => (14,13,14), 120 => (15,15,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (14,14,14), 137 => (11,11,14), 138 => (5,5,15), 139 => (0,0,3), 140 => (0,2,15), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			26 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,15), 21 => (0,0,2), 22 => (5,5,15), 23 => (11,11,14), 24 => (14,14,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (15,15,14), 44 => (14,13,14), 45 => (13,13,14), 46 => (11,10,14), 47 => (4,3,8), 48 => (3,4,15), 49 => (0,0,8), 50 => (0,0,15), 51 => (4,1,6), 52 => (15,13,4), 53 => (11,4,0), 54 => (14,9,0), 55 => (15,10,0), 56 => (13,7,0), 57 => (12,4,0), 58 => (7,0,0), 59 => (7,2,3), 60 => (4,0,2), 61 => (11,7,0), 62 => (9,4,0), 63 => (9,6,5), 64 => (11,5,0), 65 => (11,4,0), 66 => (11,4,0), 67 => (11,4,0), 68 => (10,4,0), 69 => (8,1,0), 70 => (7,5,7), 71 => (10,14,15), 72 => (10,7,4), 73 => (13,9,1), 74 => (13,8,0), 75 => (6,0,0), 76 => (13,11,0), 77 => (12,9,0), 78 => (15,15,9), 79 => (15,15,7), 80 => (0,0,14), 81 => (2,2,14), 82 => (3,3,14), 83 => (3,3,14), 84 => (1,1,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (2,2,14), 92 => (2,2,14), 93 => (2,2,14), 94 => (1,1,14), 95 => (1,1,14), 96 => (1,1,14), 97 => (2,2,14), 98 => (1,1,14), 99 => (1,1,14), 100 => (2,2,15), 101 => (0,0,12), 102 => (0,0,8), 103 => (0,0,5), 104 => (0,0,6), 105 => (0,0,0), 106 => (0,0,0), 107 => (0,2,15), 108 => (0,1,14), 109 => (0,0,14), 110 => (0,0,8), 111 => (3,4,15), 112 => (4,3,8), 113 => (11,10,14), 114 => (13,13,14), 115 => (14,13,14), 116 => (15,15,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (14,14,14), 136 => (11,11,14), 137 => (5,5,15), 138 => (0,0,2), 139 => (0,2,15), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			27 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,15), 22 => (0,0,2), 23 => (5,5,15), 24 => (11,11,14), 25 => (14,14,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (15,15,14), 48 => (14,13,14), 49 => (13,13,14), 50 => (13,13,14), 51 => (8,6,11), 52 => (14,9,0), 53 => (3,1,6), 54 => (5,6,12), 55 => (5,7,13), 56 => (7,6,7), 57 => (9,8,4), 58 => (15,10,0), 59 => (14,7,0), 60 => (11,4,0), 61 => (8,2,0), 62 => (15,8,0), 63 => (14,8,0), 64 => (14,8,0), 65 => (14,8,0), 66 => (14,8,0), 67 => (14,8,0), 68 => (13,7,0), 69 => (12,6,0), 70 => (12,6,0), 71 => (9,2,0), 72 => (13,8,0), 73 => (13,8,0), 74 => (14,9,0), 75 => (9,3,0), 76 => (9,2,0), 77 => (8,2,0), 78 => (7,0,0), 79 => (7,1,1), 80 => (3,2,10), 81 => (0,1,14), 82 => (4,4,14), 83 => (2,2,14), 84 => (1,1,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (2,2,14), 92 => (2,2,14), 93 => (1,1,14), 94 => (2,2,14), 95 => (4,4,14), 96 => (2,2,14), 97 => (1,1,14), 98 => (2,2,14), 99 => (2,2,14), 100 => (1,1,14), 101 => (1,1,14), 102 => (1,1,15), 103 => (0,0,0), 104 => (0,0,0), 105 => (0,0,0), 106 => (3,4,12), 107 => (4,4,9), 108 => (5,5,13), 109 => (13,13,14), 110 => (13,13,14), 111 => (14,13,14), 112 => (15,15,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (14,14,14), 135 => (11,11,14), 136 => (5,5,15), 137 => (0,0,2), 138 => (0,2,15), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			28 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,15), 23 => (0,0,2), 24 => (5,5,15), 25 => (11,11,14), 26 => (14,14,14), 27 => (14,14,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,15,15), 52 => (11,6,0), 53 => (10,2,0), 54 => (7,10,15), 55 => (9,11,14), 56 => (8,11,14), 57 => (8,11,15), 58 => (6,8,15), 59 => (9,7,4), 60 => (15,9,0), 61 => (14,8,0), 62 => (14,10,0), 63 => (14,8,0), 64 => (14,7,0), 65 => (14,8,0), 66 => (14,8,0), 67 => (14,8,0), 68 => (14,8,0), 69 => (14,8,0), 70 => (12,6,0), 71 => (12,6,0), 72 => (12,6,0), 73 => (8,1,0), 74 => (9,3,0), 75 => (11,5,0), 76 => (8,3,4), 77 => (8,5,8), 78 => (2,4,15), 79 => (3,3,15), 80 => (2,0,9), 81 => (8,4,4), 82 => (4,3,9), 83 => (1,1,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (2,2,14), 92 => (1,1,14), 93 => (1,1,14), 94 => (2,2,14), 95 => (3,3,14), 96 => (4,4,14), 97 => (1,1,14), 98 => (2,2,14), 99 => (1,1,14), 100 => (2,2,14), 101 => (5,5,14), 102 => (4,4,14), 103 => (0,0,15), 104 => (0,0,0), 105 => (3,3,2), 106 => (15,15,15), 107 => (15,15,14), 108 => (14,14,14), 109 => (14,14,14), 110 => (14,14,14), 111 => (14,14,14), 112 => (14,14,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (14,14,14), 133 => (14,14,14), 134 => (11,11,14), 135 => (5,5,15), 136 => (0,0,2), 137 => (0,2,15), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			29 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,15), 24 => (0,0,2), 25 => (5,5,15), 26 => (11,11,14), 27 => (13,13,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,15), 52 => (11,7,2), 53 => (12,5,0), 54 => (9,10,11), 55 => (13,14,14), 56 => (15,15,14), 57 => (6,8,12), 58 => (7,9,13), 59 => (8,9,13), 60 => (13,6,0), 61 => (14,9,0), 62 => (14,8,0), 63 => (14,7,0), 64 => (14,8,0), 65 => (14,8,0), 66 => (14,8,0), 67 => (14,8,0), 68 => (14,8,0), 69 => (14,8,0), 70 => (14,8,0), 71 => (12,6,0), 72 => (11,5,0), 73 => (14,11,0), 74 => (13,6,0), 75 => (9,2,0), 76 => (9,1,0), 77 => (8,0,0), 78 => (13,4,0), 79 => (9,14,0), 80 => (4,9,5), 81 => (2,2,15), 82 => (1,1,14), 83 => (2,2,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (2,2,14), 91 => (0,0,14), 92 => (5,5,11), 93 => (8,8,5), 94 => (4,4,6), 95 => (0,0,10), 96 => (2,2,14), 97 => (3,3,14), 98 => (1,1,14), 99 => (1,1,14), 100 => (5,5,14), 101 => (11,11,14), 102 => (7,7,14), 103 => (1,1,14), 104 => (1,1,11), 105 => (2,2,9), 106 => (6,6,13), 107 => (15,15,14), 108 => (15,15,14), 109 => (14,14,14), 110 => (14,14,14), 111 => (14,14,14), 112 => (14,14,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (13,13,14), 133 => (11,11,14), 134 => (5,5,15), 135 => (0,0,2), 136 => (0,2,15), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			30 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,15), 25 => (0,0,2), 26 => (5,5,15), 27 => (9,9,14), 28 => (13,13,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (11,8,6), 53 => (15,10,0), 54 => (8,3,2), 55 => (13,15,15), 56 => (10,11,14), 57 => (9,12,14), 58 => (12,14,15), 59 => (11,4,0), 60 => (14,11,4), 61 => (14,10,1), 62 => (14,8,0), 63 => (14,7,0), 64 => (14,8,0), 65 => (14,8,0), 66 => (14,8,0), 67 => (14,8,0), 68 => (14,8,0), 69 => (14,8,0), 70 => (14,8,0), 71 => (13,7,0), 72 => (11,5,0), 73 => (7,0,0), 74 => (5,5,0), 75 => (7,15,0), 76 => (7,15,0), 77 => (8,15,0), 78 => (6,6,0), 79 => (9,0,0), 80 => (2,0,10), 81 => (2,2,15), 82 => (1,1,14), 83 => (2,2,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (2,2,14), 90 => (0,0,14), 91 => (8,8,9), 92 => (14,14,13), 93 => (14,14,14), 94 => (15,15,15), 95 => (11,11,8), 96 => (0,0,10), 97 => (2,2,14), 98 => (1,1,14), 99 => (1,1,14), 100 => (3,3,14), 101 => (7,7,14), 102 => (5,5,14), 103 => (1,1,14), 104 => (1,1,13), 105 => (3,3,14), 106 => (4,4,14), 107 => (1,1,13), 108 => (0,0,12), 109 => (6,6,12), 110 => (11,11,13), 111 => (15,15,14), 112 => (14,14,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (13,13,14), 132 => (9,9,14), 133 => (5,5,15), 134 => (0,0,2), 135 => (0,2,15), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			31 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,15), 26 => (0,0,3), 27 => (0,0,8), 28 => (10,10,15), 29 => (11,11,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (8,9,15), 53 => (12,7,0), 54 => (9,1,0), 55 => (12,15,15), 56 => (9,11,14), 57 => (14,14,14), 58 => (10,7,6), 59 => (13,9,2), 60 => (14,15,15), 61 => (14,11,6), 62 => (14,8,0), 63 => (14,7,0), 64 => (14,8,0), 65 => (14,7,0), 66 => (14,7,0), 67 => (14,8,0), 68 => (14,8,0), 69 => (14,8,0), 70 => (14,8,0), 71 => (13,7,0), 72 => (12,6,0), 73 => (10,7,0), 74 => (7,15,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,15,0), 80 => (4,0,5), 81 => (4,2,10), 82 => (1,1,14), 83 => (2,2,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (2,2,14), 89 => (1,1,14), 90 => (5,5,11), 91 => (14,14,13), 92 => (14,14,14), 93 => (14,14,14), 94 => (14,14,14), 95 => (15,15,15), 96 => (9,9,7), 97 => (0,0,13), 98 => (2,2,14), 99 => (2,2,14), 100 => (1,1,14), 101 => (2,2,14), 102 => (2,2,14), 103 => (1,1,14), 104 => (0,0,12), 105 => (0,0,13), 106 => (1,1,14), 107 => (1,1,14), 108 => (3,3,14), 109 => (2,2,14), 110 => (1,1,13), 111 => (2,2,12), 112 => (15,15,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (11,11,14), 131 => (10,10,15), 132 => (0,0,8), 133 => (0,0,3), 134 => (0,2,15), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			32 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,15), 27 => (0,1,9), 28 => (0,0,8), 29 => (5,5,14), 30 => (10,10,14), 31 => (13,13,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (4,4,14), 53 => (7,4,7), 54 => (15,10,0), 55 => (5,3,7), 56 => (11,13,15), 57 => (9,13,15), 58 => (11,3,0), 59 => (14,11,4), 60 => (14,11,6), 61 => (14,10,1), 62 => (14,8,0), 63 => (14,7,0), 64 => (14,8,0), 65 => (12,7,2), 66 => (10,9,7), 67 => (11,7,3), 68 => (14,8,0), 69 => (14,7,0), 70 => (13,8,1), 71 => (11,10,8), 72 => (14,7,0), 73 => (11,3,0), 74 => (7,15,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,15,0), 80 => (0,0,15), 81 => (5,3,7), 82 => (4,2,9), 83 => (1,1,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (1,1,14), 89 => (2,2,12), 90 => (14,14,12), 91 => (14,14,14), 92 => (10,10,10), 93 => (11,11,11), 94 => (14,14,14), 95 => (14,14,14), 96 => (12,12,12), 97 => (3,3,8), 98 => (1,1,14), 99 => (2,2,14), 100 => (2,2,14), 101 => (1,1,14), 102 => (3,3,14), 103 => (2,2,14), 104 => (1,1,14), 105 => (1,1,10), 106 => (3,3,9), 107 => (2,2,12), 108 => (1,1,14), 109 => (1,1,14), 110 => (2,2,14), 111 => (3,3,14), 112 => (0,0,13), 113 => (10,10,13), 114 => (15,15,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (13,13,14), 129 => (10,10,14), 130 => (5,5,14), 131 => (0,0,8), 132 => (0,1,9), 133 => (0,2,15), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			33 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,1,14), 26 => (0,1,14), 27 => (0,2,14), 28 => (0,1,10), 29 => (0,0,3), 30 => (2,1,14), 31 => (9,9,14), 32 => (11,11,14), 33 => (13,13,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (9,9,14), 52 => (4,4,14), 53 => (4,5,15), 54 => (11,5,0), 55 => (12,6,0), 56 => (8,9,12), 57 => (9,7,7), 58 => (13,6,0), 59 => (14,11,5), 60 => (14,10,1), 61 => (14,8,0), 62 => (14,7,0), 63 => (14,8,0), 64 => (12,5,0), 65 => (12,15,15), 66 => (13,14,15), 67 => (11,11,11), 68 => (13,6,0), 69 => (14,8,0), 70 => (12,8,4), 71 => (12,15,15), 72 => (12,5,0), 73 => (11,3,0), 74 => (7,15,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,15,0), 80 => (0,0,15), 81 => (9,9,6), 82 => (3,3,14), 83 => (1,1,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (2,2,14), 88 => (0,0,13), 89 => (8,8,10), 90 => (14,14,14), 91 => (14,14,14), 92 => (4,4,4), 93 => (0,0,0), 94 => (13,13,13), 95 => (14,14,14), 96 => (15,15,14), 97 => (4,4,10), 98 => (1,1,14), 99 => (2,2,14), 100 => (2,2,14), 101 => (1,1,14), 102 => (1,1,14), 103 => (1,1,14), 104 => (2,2,13), 105 => (8,8,6), 106 => (12,12,11), 107 => (9,9,7), 108 => (5,5,7), 109 => (1,1,15), 110 => (1,1,14), 111 => (0,0,15), 112 => (3,3,8), 113 => (10,10,9), 114 => (6,6,6), 115 => (12,12,12), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (13,13,14), 127 => (11,11,14), 128 => (9,9,14), 129 => (2,1,14), 130 => (0,0,3), 131 => (0,1,10), 132 => (0,2,14), 133 => (0,1,14), 134 => (0,1,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			34 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (1,1,8), 25 => (4,4,8), 26 => (5,6,14), 27 => (0,1,13), 28 => (0,0,9), 29 => (0,1,15), 30 => (0,0,4), 31 => (0,0,8), 32 => (5,5,14), 33 => (9,9,14), 34 => (11,11,14), 35 => (13,13,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (4,4,14), 52 => (7,7,15), 53 => (3,1,5), 54 => (11,8,0), 55 => (14,7,0), 56 => (7,3,3), 57 => (11,4,0), 58 => (12,6,0), 59 => (14,9,0), 60 => (14,8,0), 61 => (14,7,0), 62 => (14,8,0), 63 => (14,8,0), 64 => (13,10,8), 65 => (13,14,14), 66 => (14,14,14), 67 => (14,15,15), 68 => (13,7,0), 69 => (14,8,0), 70 => (4,1,0), 71 => (10,11,15), 72 => (12,5,0), 73 => (11,3,0), 74 => (7,15,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,15,0), 80 => (1,2,11), 81 => (8,8,7), 82 => (8,8,10), 83 => (0,0,14), 84 => (2,2,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (1,1,14), 88 => (1,1,11), 89 => (14,14,13), 90 => (14,14,14), 91 => (14,14,14), 92 => (13,13,13), 93 => (3,3,3), 94 => (8,8,8), 95 => (14,14,14), 96 => (15,15,14), 97 => (4,4,10), 98 => (1,1,14), 99 => (2,2,14), 100 => (2,2,14), 101 => (1,1,14), 102 => (7,7,9), 103 => (9,9,7), 104 => (9,9,8), 105 => (15,15,15), 106 => (14,14,14), 107 => (13,13,13), 108 => (8,8,7), 109 => (4,4,6), 110 => (1,1,13), 111 => (6,6,8), 112 => (15,15,14), 113 => (11,11,11), 114 => (8,8,8), 115 => (9,9,9), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (13,13,14), 125 => (11,11,14), 126 => (9,9,14), 127 => (5,5,14), 128 => (0,0,8), 129 => (0,0,4), 130 => (0,1,15), 131 => (0,0,9), 132 => (0,1,13), 133 => (5,6,14), 134 => (4,4,8), 135 => (1,1,8), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			35 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,0,3), 25 => (6,6,15), 26 => (12,12,14), 27 => (13,13,14), 28 => (13,13,14), 29 => (5,5,13), 30 => (4,5,10), 31 => (3,4,10), 32 => (0,0,3), 33 => (0,0,8), 34 => (4,4,14), 35 => (8,8,14), 36 => (10,10,14), 37 => (13,13,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (9,9,14), 51 => (5,5,14), 52 => (1,2,15), 53 => (12,7,0), 54 => (8,7,4), 55 => (10,7,3), 56 => (14,7,0), 57 => (12,6,0), 58 => (11,5,0), 59 => (14,8,0), 60 => (14,7,0), 61 => (14,8,0), 62 => (14,8,0), 63 => (12,5,0), 64 => (2,0,3), 65 => (15,15,15), 66 => (14,14,14), 67 => (14,14,15), 68 => (14,9,3), 69 => (14,7,0), 70 => (15,13,9), 71 => (5,6,7), 72 => (12,5,0), 73 => (10,6,0), 74 => (7,14,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (4,7,7), 81 => (5,4,11), 82 => (15,15,13), 83 => (8,8,9), 84 => (0,0,14), 85 => (2,2,14), 86 => (2,2,14), 87 => (0,0,13), 88 => (8,8,10), 89 => (14,14,14), 90 => (14,14,14), 91 => (14,14,14), 92 => (8,8,8), 93 => (0,0,0), 94 => (0,0,0), 95 => (15,15,15), 96 => (15,15,14), 97 => (3,3,10), 98 => (0,0,15), 99 => (0,1,14), 100 => (1,1,15), 101 => (0,0,15), 102 => (12,12,10), 103 => (14,14,14), 104 => (8,8,8), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (10,10,10), 109 => (7,7,6), 110 => (8,8,7), 111 => (13,13,13), 112 => (9,9,9), 113 => (8,8,8), 114 => (2,2,2), 115 => (5,5,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (13,13,14), 123 => (10,10,14), 124 => (8,8,14), 125 => (4,4,14), 126 => (0,0,8), 127 => (0,0,3), 128 => (3,4,10), 129 => (4,5,10), 130 => (5,5,13), 131 => (13,13,14), 132 => (13,13,14), 133 => (12,12,14), 134 => (6,6,15), 135 => (0,0,3), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			36 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,1,10), 25 => (0,0,8), 26 => (9,9,14), 27 => (13,13,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (15,15,14), 31 => (14,13,14), 32 => (13,13,15), 33 => (9,9,9), 34 => (5,5,8), 35 => (7,7,13), 36 => (10,10,14), 37 => (11,11,14), 38 => (12,12,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (14,13,14), 50 => (4,4,14), 51 => (6,6,15), 52 => (3,1,5), 53 => (14,12,0), 54 => (11,11,0), 55 => (1,2,15), 56 => (11,4,0), 57 => (12,6,0), 58 => (11,5,0), 59 => (12,6,0), 60 => (14,8,0), 61 => (14,8,0), 62 => (14,8,0), 63 => (12,5,0), 64 => (10,12,15), 65 => (10,12,14), 66 => (14,14,14), 67 => (14,14,15), 68 => (14,9,3), 69 => (14,8,0), 70 => (5,2,0), 71 => (6,7,8), 72 => (13,5,0), 73 => (8,9,0), 74 => (7,14,0), 75 => (8,14,0), 76 => (8,14,0), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,15,0), 81 => (2,3,12), 82 => (11,11,13), 83 => (14,14,13), 84 => (8,8,9), 85 => (1,1,15), 86 => (1,1,14), 87 => (1,1,11), 88 => (14,14,13), 89 => (14,14,14), 90 => (14,14,14), 91 => (14,14,14), 92 => (5,5,5), 93 => (0,0,0), 94 => (0,0,0), 95 => (15,15,15), 96 => (14,15,14), 97 => (7,6,9), 98 => (14,11,7), 99 => (14,11,8), 100 => (10,5,1), 101 => (5,4,6), 102 => (15,15,15), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (12,12,12), 109 => (8,8,8), 110 => (5,5,5), 111 => (10,10,10), 112 => (7,7,7), 113 => (7,7,7), 114 => (15,15,15), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (12,12,14), 122 => (11,11,14), 123 => (10,10,14), 124 => (7,7,13), 125 => (5,5,8), 126 => (9,9,9), 127 => (13,13,15), 128 => (14,13,14), 129 => (15,15,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (13,13,14), 133 => (9,9,14), 134 => (0,0,8), 135 => (0,1,10), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			37 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,15), 25 => (0,0,3), 26 => (5,5,15), 27 => (11,11,14), 28 => (14,14,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (15,15,14), 42 => (10,12,14), 43 => (8,10,14), 44 => (8,10,14), 45 => (7,10,14), 46 => (8,11,14), 47 => (7,10,14), 48 => (10,11,14), 49 => (9,11,14), 50 => (4,4,14), 51 => (1,1,14), 52 => (12,6,0), 53 => (14,15,0), 54 => (11,11,10), 55 => (3,3,2), 56 => (12,7,0), 57 => (12,5,0), 58 => (11,5,0), 59 => (12,6,0), 60 => (14,8,0), 61 => (14,8,0), 62 => (14,8,0), 63 => (12,5,0), 64 => (7,8,11), 65 => (7,7,8), 66 => (14,14,14), 67 => (14,14,15), 68 => (14,9,3), 69 => (14,8,0), 70 => (7,4,2), 71 => (5,6,7), 72 => (12,4,0), 73 => (8,8,0), 74 => (8,13,3), 75 => (2,5,0), 76 => (7,9,6), 77 => (8,13,4), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,14,0), 81 => (7,12,2), 82 => (4,3,15), 83 => (15,15,14), 84 => (14,14,13), 85 => (1,1,3), 86 => (4,4,10), 87 => (8,8,10), 88 => (14,14,14), 89 => (14,14,14), 90 => (14,14,14), 91 => (14,14,14), 92 => (15,15,15), 93 => (0,0,0), 94 => (0,0,0), 95 => (15,15,15), 96 => (13,12,12), 97 => (14,9,6), 98 => (14,11,10), 99 => (14,11,10), 100 => (15,10,7), 101 => (10,11,11), 102 => (14,14,14), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (14,14,14), 109 => (9,9,9), 110 => (8,8,8), 111 => (10,10,10), 112 => (7,7,7), 113 => (15,15,15), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (14,14,14), 132 => (11,11,14), 133 => (5,5,15), 134 => (0,0,3), 135 => (0,2,15), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			38 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,15), 26 => (0,0,2), 27 => (8,8,15), 28 => (12,12,14), 29 => (14,14,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (13,13,14), 41 => (4,5,11), 42 => (6,7,11), 43 => (8,10,14), 44 => (11,13,14), 45 => (14,14,14), 46 => (14,14,14), 47 => (13,14,14), 48 => (11,13,14), 49 => (11,13,14), 50 => (9,11,14), 51 => (3,5,15), 52 => (14,11,0), 53 => (14,14,0), 54 => (9,9,0), 55 => (15,15,0), 56 => (13,12,0), 57 => (11,4,0), 58 => (12,5,0), 59 => (12,5,0), 60 => (12,5,0), 61 => (13,7,0), 62 => (14,8,0), 63 => (12,6,0), 64 => (0,0,1), 65 => (6,6,5), 66 => (14,14,14), 67 => (14,14,15), 68 => (14,9,2), 69 => (14,6,0), 70 => (9,8,6), 71 => (10,13,15), 72 => (9,12,15), 73 => (11,13,15), 74 => (2,1,4), 75 => (0,0,2), 76 => (7,6,8), 77 => (5,9,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,14,0), 81 => (8,15,0), 82 => (3,6,7), 83 => (13,12,15), 84 => (15,15,15), 85 => (4,4,4), 86 => (6,6,6), 87 => (15,15,15), 88 => (14,14,14), 89 => (14,14,14), 90 => (14,14,14), 91 => (14,14,14), 92 => (14,14,14), 93 => (14,14,14), 94 => (9,10,10), 95 => (13,14,14), 96 => (12,7,5), 97 => (14,10,8), 98 => (14,9,7), 99 => (10,5,3), 100 => (10,8,7), 101 => (14,15,15), 102 => (14,14,14), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (14,14,14), 109 => (9,9,9), 110 => (10,10,10), 111 => (9,9,9), 112 => (9,9,9), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,14,14), 131 => (12,12,14), 132 => (8,8,15), 133 => (0,0,2), 134 => (0,2,15), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			39 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,1,10), 27 => (0,0,8), 28 => (9,9,14), 29 => (13,13,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (8,9,12), 41 => (15,15,14), 42 => (15,14,14), 43 => (12,12,12), 44 => (6,7,11), 45 => (11,13,14), 46 => (14,14,14), 47 => (14,14,14), 48 => (14,14,14), 49 => (13,14,14), 50 => (13,14,14), 51 => (10,13,14), 52 => (8,10,12), 53 => (15,14,0), 54 => (14,14,0), 55 => (14,14,0), 56 => (12,13,4), 57 => (7,5,9), 58 => (10,8,7), 59 => (6,6,8), 60 => (6,10,15), 61 => (10,8,6), 62 => (10,9,7), 63 => (15,8,0), 64 => (0,0,3), 65 => (13,13,14), 66 => (14,14,14), 67 => (14,14,14), 68 => (13,13,13), 69 => (14,14,15), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (12,14,14), 74 => (9,12,15), 75 => (7,9,14), 76 => (5,5,12), 77 => (8,15,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,14,0), 81 => (8,14,0), 82 => (9,15,0), 83 => (3,4,10), 84 => (15,15,14), 85 => (11,11,11), 86 => (3,3,3), 87 => (14,13,13), 88 => (14,14,14), 89 => (14,14,14), 90 => (14,14,14), 91 => (14,14,14), 92 => (14,14,14), 93 => (14,14,14), 94 => (13,13,13), 95 => (12,9,7), 96 => (14,10,8), 97 => (14,10,8), 98 => (9,5,3), 99 => (14,10,8), 100 => (10,8,7), 101 => (13,13,13), 102 => (14,14,14), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (14,14,14), 109 => (9,9,9), 110 => (9,9,9), 111 => (5,5,5), 112 => (15,15,15), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (13,13,14), 131 => (9,9,14), 132 => (0,0,8), 133 => (0,1,10), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			40 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,15), 27 => (0,0,3), 28 => (5,5,15), 29 => (11,11,14), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (15,15,14), 45 => (6,7,11), 46 => (10,13,14), 47 => (13,14,14), 48 => (14,14,14), 49 => (14,14,14), 50 => (13,14,14), 51 => (11,14,14), 52 => (11,13,14), 53 => (8,10,12), 54 => (14,14,0), 55 => (14,14,0), 56 => (14,14,0), 57 => (14,12,0), 58 => (6,5,8), 59 => (12,13,15), 60 => (9,10,12), 61 => (14,15,15), 62 => (14,14,14), 63 => (10,13,15), 64 => (12,15,15), 65 => (13,14,14), 66 => (14,14,14), 67 => (14,14,14), 68 => (14,14,15), 69 => (14,14,14), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (13,14,14), 74 => (11,13,14), 75 => (8,11,14), 76 => (8,8,14), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,14,0), 81 => (8,14,0), 82 => (5,8,1), 83 => (3,7,0), 84 => (0,0,5), 85 => (8,8,8), 86 => (0,1,1), 87 => (10,7,5), 88 => (13,9,8), 89 => (12,10,9), 90 => (12,13,13), 91 => (14,14,15), 92 => (14,15,15), 93 => (12,10,9), 94 => (13,8,6), 95 => (14,10,8), 96 => (14,10,8), 97 => (9,5,3), 98 => (12,8,6), 99 => (14,10,8), 100 => (11,9,8), 101 => (10,11,10), 102 => (14,14,14), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (14,14,14), 108 => (12,12,12), 109 => (9,9,9), 110 => (8,8,8), 111 => (8,8,10), 112 => (14,14,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (11,11,14), 131 => (5,5,15), 132 => (0,0,3), 133 => (0,2,15), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			41 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,15), 28 => (0,0,3), 29 => (5,5,14), 30 => (11,11,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (6,8,12), 45 => (11,11,13), 46 => (8,10,14), 47 => (11,13,14), 48 => (13,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (13,14,14), 53 => (10,12,15), 54 => (10,11,7), 55 => (14,14,0), 56 => (14,14,0), 57 => (10,12,8), 58 => (10,8,9), 59 => (13,14,14), 60 => (14,14,14), 61 => (14,14,14), 62 => (14,14,14), 63 => (14,14,14), 64 => (14,14,14), 65 => (14,14,14), 66 => (13,14,14), 67 => (14,13,11), 68 => (9,7,6), 69 => (7,10,10), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (12,14,14), 74 => (11,13,14), 75 => (10,12,15), 76 => (6,8,4), 77 => (8,14,0), 78 => (8,14,0), 79 => (8,14,0), 80 => (8,14,0), 81 => (8,15,0), 82 => (0,0,2), 83 => (8,8,8), 84 => (7,7,7), 85 => (0,0,0), 86 => (0,0,0), 87 => (13,8,6), 88 => (14,10,8), 89 => (14,10,7), 90 => (12,8,6), 91 => (12,8,6), 92 => (12,8,5), 93 => (14,10,7), 94 => (14,10,8), 95 => (14,10,8), 96 => (11,7,5), 97 => (13,9,7), 98 => (14,10,8), 99 => (15,11,8), 100 => (7,3,4), 101 => (5,5,9), 102 => (15,15,14), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (14,14,14), 107 => (13,13,13), 108 => (9,9,9), 109 => (10,10,10), 110 => (7,7,7), 111 => (7,7,9), 112 => (14,14,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (11,11,14), 130 => (5,5,14), 131 => (0,0,3), 132 => (0,2,15), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			42 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,1,10), 29 => (0,0,8), 30 => (8,8,15), 31 => (11,11,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (15,14,14), 45 => (8,9,12), 46 => (8,9,12), 47 => (10,12,14), 48 => (12,14,14), 49 => (14,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (14,14,14), 53 => (12,14,14), 54 => (7,10,15), 55 => (13,13,1), 56 => (10,11,8), 57 => (10,11,11), 58 => (5,6,12), 59 => (11,13,14), 60 => (14,14,14), 61 => (14,14,14), 62 => (14,14,14), 63 => (14,14,14), 64 => (14,14,14), 65 => (14,14,14), 66 => (14,15,15), 67 => (6,0,0), 68 => (9,1,0), 69 => (7,5,6), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (11,14,14), 74 => (8,9,14), 75 => (5,5,7), 76 => (8,15,0), 77 => (8,14,0), 78 => (7,14,0), 79 => (7,14,0), 80 => (8,14,0), 81 => (8,14,0), 82 => (6,11,0), 83 => (3,1,4), 84 => (1,0,2), 85 => (4,6,3), 86 => (6,3,3), 87 => (13,8,6), 88 => (13,9,7), 89 => (14,10,8), 90 => (14,10,8), 91 => (14,10,8), 92 => (14,10,8), 93 => (14,10,8), 94 => (14,10,8), 95 => (14,10,8), 96 => (14,10,8), 97 => (14,10,8), 98 => (15,11,9), 99 => (7,4,4), 100 => (0,0,14), 101 => (3,3,9), 102 => (11,11,10), 103 => (14,14,14), 104 => (14,14,14), 105 => (14,14,14), 106 => (12,12,12), 107 => (9,9,9), 108 => (10,10,10), 109 => (9,9,9), 110 => (6,6,6), 111 => (3,3,12), 112 => (13,13,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (11,11,14), 129 => (8,8,15), 130 => (0,0,8), 131 => (0,1,10), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			43 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,1,9), 30 => (0,0,8), 31 => (8,8,15), 32 => (11,11,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,14,14), 45 => (12,11,12), 46 => (8,10,13), 47 => (10,12,14), 48 => (11,13,14), 49 => (13,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (14,14,14), 53 => (13,14,14), 54 => (10,13,14), 55 => (9,10,11), 56 => (15,15,0), 57 => (7,7,6), 58 => (6,7,12), 59 => (8,9,11), 60 => (14,14,14), 61 => (14,14,14), 62 => (14,14,14), 63 => (14,14,14), 64 => (14,14,14), 65 => (14,14,14), 66 => (14,14,14), 67 => (12,13,15), 68 => (7,2,0), 69 => (12,8,5), 70 => (14,14,14), 71 => (14,14,14), 72 => (10,11,14), 73 => (6,7,9), 74 => (7,12,1), 75 => (8,15,0), 76 => (8,14,0), 77 => (6,11,0), 78 => (9,8,14), 79 => (10,8,14), 80 => (6,11,0), 81 => (8,14,0), 82 => (8,14,0), 83 => (8,15,0), 84 => (8,15,0), 85 => (8,15,0), 86 => (6,11,0), 87 => (7,5,1), 88 => (12,7,6), 89 => (12,8,6), 90 => (13,9,7), 91 => (14,10,8), 92 => (14,10,8), 93 => (14,10,8), 94 => (14,10,8), 95 => (14,10,8), 96 => (15,11,9), 97 => (14,9,7), 98 => (2,0,0), 99 => (0,0,5), 100 => (0,0,8), 101 => (0,0,12), 102 => (5,5,7), 103 => (10,10,10), 104 => (12,12,12), 105 => (10,10,10), 106 => (9,9,9), 107 => (10,10,10), 108 => (9,9,9), 109 => (7,7,7), 110 => (6,6,5), 111 => (3,3,7), 112 => (12,12,14), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (11,11,14), 128 => (8,8,15), 129 => (0,0,8), 130 => (0,1,9), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			44 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,1,9), 31 => (0,0,8), 32 => (8,8,15), 33 => (11,11,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (15,15,14), 42 => (9,8,11), 43 => (9,9,11), 44 => (9,8,11), 45 => (15,15,14), 46 => (5,6,11), 47 => (8,11,14), 48 => (10,12,14), 49 => (11,14,14), 50 => (14,14,14), 51 => (14,14,14), 52 => (14,14,14), 53 => (14,14,14), 54 => (12,13,14), 55 => (8,10,15), 56 => (13,14,0), 57 => (6,6,15), 58 => (5,5,14), 59 => (11,13,14), 60 => (14,14,14), 61 => (13,14,14), 62 => (11,14,14), 63 => (12,14,14), 64 => (13,14,14), 65 => (13,14,14), 66 => (14,14,14), 67 => (14,14,14), 68 => (13,14,15), 69 => (14,15,15), 70 => (15,14,14), 71 => (9,10,15), 72 => (6,11,0), 73 => (8,14,0), 74 => (8,14,0), 75 => (8,14,0), 76 => (6,12,0), 77 => (12,11,15), 78 => (13,14,14), 79 => (13,14,14), 80 => (12,11,15), 81 => (6,11,0), 82 => (8,14,0), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,15,0), 88 => (7,8,0), 89 => (8,6,2), 90 => (9,4,3), 91 => (13,8,7), 92 => (14,9,7), 93 => (14,9,7), 94 => (13,8,6), 95 => (10,6,4), 96 => (4,1,0), 97 => (1,0,0), 98 => (0,0,7), 99 => (0,0,14), 100 => (2,2,14), 101 => (1,1,13), 102 => (0,0,13), 103 => (4,4,3), 104 => (8,8,8), 105 => (9,9,9), 106 => (9,9,9), 107 => (9,9,9), 108 => (7,7,7), 109 => (6,6,6), 110 => (9,9,9), 111 => (7,7,5), 112 => (6,6,13), 113 => (14,14,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (11,11,14), 127 => (8,8,15), 128 => (0,0,8), 129 => (0,1,9), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			45 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,1,9), 32 => (0,0,8), 33 => (8,8,15), 34 => (11,11,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (12,12,12), 41 => (6,7,11), 42 => (10,12,14), 43 => (10,12,14), 44 => (10,12,14), 45 => (6,7,11), 46 => (6,6,10), 47 => (9,11,14), 48 => (9,11,14), 49 => (12,14,14), 50 => (13,14,14), 51 => (14,14,14), 52 => (14,14,14), 53 => (14,14,14), 54 => (13,14,14), 55 => (10,12,14), 56 => (10,11,10), 57 => (5,4,14), 58 => (10,12,14), 59 => (7,8,11), 60 => (13,14,14), 61 => (11,14,14), 62 => (8,10,14), 63 => (7,8,13), 64 => (8,9,13), 65 => (11,13,15), 66 => (12,14,15), 67 => (15,15,15), 68 => (14,15,15), 69 => (11,12,14), 70 => (6,9,9), 71 => (7,12,1), 72 => (8,14,0), 73 => (8,14,0), 74 => (8,14,0), 75 => (8,14,0), 76 => (8,6,13), 77 => (6,6,10), 78 => (10,13,14), 79 => (14,14,14), 80 => (14,14,14), 81 => (8,9,15), 82 => (7,11,1), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,14,0), 88 => (8,14,0), 89 => (7,14,0), 90 => (7,15,0), 91 => (8,9,0), 92 => (2,0,0), 93 => (1,0,0), 94 => (1,0,0), 95 => (0,0,0), 96 => (5,2,0), 97 => (3,1,9), 98 => (5,2,7), 99 => (0,1,15), 100 => (1,1,14), 101 => (1,1,15), 102 => (4,2,6), 103 => (7,7,7), 104 => (10,10,10), 105 => (11,11,11), 106 => (10,10,10), 107 => (11,11,11), 108 => (9,9,9), 109 => (12,12,12), 110 => (9,9,8), 111 => (5,5,6), 112 => (0,0,13), 113 => (15,15,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (11,11,14), 126 => (8,8,15), 127 => (0,0,8), 128 => (0,1,9), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			46 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,1,10), 33 => (0,0,2), 34 => (5,5,15), 35 => (10,10,14), 36 => (13,13,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (12,12,12), 40 => (6,8,13), 41 => (9,11,14), 42 => (8,10,14), 43 => (8,10,14), 44 => (10,12,14), 45 => (10,13,14), 46 => (5,4,8), 47 => (8,10,14), 48 => (10,12,14), 49 => (11,13,14), 50 => (11,14,14), 51 => (14,14,14), 52 => (14,14,14), 53 => (14,14,14), 54 => (12,13,14), 55 => (10,12,14), 56 => (8,9,14), 57 => (5,7,14), 58 => (4,4,10), 59 => (12,15,9), 60 => (10,12,15), 61 => (6,6,10), 62 => (8,2,0), 63 => (10,4,0), 64 => (4,0,0), 65 => (0,1,4), 66 => (1,1,3), 67 => (0,1,3), 68 => (5,1,3), 69 => (5,1,3), 70 => (5,0,0), 71 => (7,11,0), 72 => (8,13,4), 73 => (8,14,0), 74 => (7,14,0), 75 => (7,13,2), 76 => (7,8,13), 77 => (15,15,15), 78 => (11,11,12), 79 => (11,13,14), 80 => (14,14,14), 81 => (13,13,15), 82 => (6,8,4), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,14,0), 88 => (8,14,0), 89 => (8,14,0), 90 => (8,15,0), 91 => (4,3,0), 92 => (4,2,0), 93 => (5,2,0), 94 => (9,5,3), 95 => (10,6,4), 96 => (13,8,6), 97 => (12,8,5), 98 => (13,9,5), 99 => (9,5,5), 100 => (1,1,12), 101 => (4,2,7), 102 => (15,10,6), 103 => (10,11,11), 104 => (9,9,9), 105 => (14,14,14), 106 => (15,15,15), 107 => (15,15,15), 108 => (12,12,12), 109 => (8,8,8), 110 => (5,5,8), 111 => (0,0,12), 112 => (1,1,13), 113 => (6,6,12), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (13,13,14), 124 => (10,10,14), 125 => (5,5,15), 126 => (0,0,2), 127 => (0,1,10), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			47 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,15), 34 => (0,0,2), 35 => (2,1,14), 36 => (9,9,14), 37 => (11,11,14), 38 => (15,15,14), 39 => (9,9,11), 40 => (9,9,11), 41 => (10,9,11), 42 => (5,6,11), 43 => (7,10,14), 44 => (8,10,14), 45 => (10,13,14), 46 => (5,4,9), 47 => (8,10,14), 48 => (8,10,14), 49 => (11,13,14), 50 => (12,14,14), 51 => (13,14,14), 52 => (14,14,14), 53 => (14,14,14), 54 => (11,13,14), 55 => (10,10,10), 56 => (7,10,15), 57 => (3,4,12), 58 => (6,6,14), 59 => (10,11,15), 60 => (6,9,9), 61 => (8,0,0), 62 => (14,9,0), 63 => (14,13,11), 64 => (14,10,1), 65 => (9,4,1), 66 => (6,6,10), 67 => (5,1,2), 68 => (6,8,13), 69 => (6,8,13), 70 => (5,0,2), 71 => (6,9,15), 72 => (6,3,1), 73 => (7,13,2), 74 => (8,12,7), 75 => (8,11,12), 76 => (5,7,5), 77 => (7,9,12), 78 => (6,6,10), 79 => (11,13,14), 80 => (13,13,14), 81 => (10,12,15), 82 => (6,9,4), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,14,0), 88 => (8,14,0), 89 => (8,15,0), 90 => (5,7,0), 91 => (7,2,1), 92 => (7,3,1), 93 => (11,7,5), 94 => (12,8,6), 95 => (12,8,6), 96 => (11,7,5), 97 => (12,8,6), 98 => (14,11,9), 99 => (14,13,11), 100 => (13,8,4), 101 => (2,0,3), 102 => (12,7,5), 103 => (12,8,6), 104 => (5,6,7), 105 => (9,9,9), 106 => (8,9,9), 107 => (8,9,9), 108 => (9,9,10), 109 => (5,5,4), 110 => (1,0,0), 111 => (0,0,13), 112 => (0,0,13), 113 => (0,0,13), 114 => (15,15,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (15,15,14), 122 => (11,11,14), 123 => (9,9,14), 124 => (2,1,14), 125 => (0,0,2), 126 => (0,2,15), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			48 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,1,14), 33 => (0,1,14), 34 => (0,2,15), 35 => (0,0,4), 36 => (0,0,8), 37 => (5,5,14), 38 => (9,9,14), 39 => (9,9,11), 40 => (15,15,14), 41 => (14,14,14), 42 => (15,15,14), 43 => (6,6,9), 44 => (6,7,11), 45 => (8,10,15), 46 => (5,5,9), 47 => (6,7,11), 48 => (7,9,14), 49 => (10,12,14), 50 => (10,13,14), 51 => (11,11,10), 52 => (14,14,14), 53 => (13,13,14), 54 => (11,13,15), 55 => (15,9,0), 56 => (10,6,3), 57 => (9,3,1), 58 => (7,8,15), 59 => (7,13,0), 60 => (6,6,0), 61 => (12,6,0), 62 => (13,7,0), 63 => (14,11,5), 64 => (14,10,0), 65 => (14,8,0), 66 => (10,5,2), 67 => (9,13,15), 68 => (9,12,14), 69 => (10,12,14), 70 => (11,14,15), 71 => (15,14,14), 72 => (11,12,15), 73 => (11,12,15), 74 => (12,11,14), 75 => (6,10,4), 76 => (7,9,8), 77 => (5,4,9), 78 => (5,5,9), 79 => (9,11,13), 80 => (10,13,15), 81 => (6,5,12), 82 => (7,12,1), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,14,0), 88 => (8,14,0), 89 => (5,11,0), 90 => (5,1,1), 91 => (7,3,1), 92 => (11,7,5), 93 => (12,8,6), 94 => (12,8,6), 95 => (12,8,6), 96 => (11,7,5), 97 => (13,9,6), 98 => (14,15,15), 99 => (14,14,15), 100 => (14,13,12), 101 => (8,4,1), 102 => (6,3,1), 103 => (13,8,6), 104 => (15,10,8), 105 => (2,2,1), 106 => (4,3,2), 107 => (4,3,2), 108 => (3,0,0), 109 => (7,3,0), 110 => (1,0,7), 111 => (3,3,5), 112 => (0,0,4), 113 => (0,0,9), 114 => (5,5,13), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (13,13,14), 121 => (9,9,14), 122 => (5,5,14), 123 => (0,0,8), 124 => (0,0,4), 125 => (0,2,15), 126 => (0,1,14), 127 => (0,1,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			49 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,1,14), 32 => (1,2,14), 33 => (6,7,14), 34 => (0,1,13), 35 => (0,0,10), 36 => (0,0,10), 37 => (0,0,4), 38 => (0,0,9), 39 => (9,9,15), 40 => (11,11,14), 41 => (13,13,14), 42 => (14,14,14), 43 => (12,12,13), 44 => (4,4,9), 45 => (6,7,11), 46 => (5,5,9), 47 => (6,6,11), 48 => (7,10,14), 49 => (8,10,14), 50 => (10,13,15), 51 => (15,7,0), 52 => (9,12,15), 53 => (12,13,14), 54 => (10,11,11), 55 => (14,10,0), 56 => (14,7,0), 57 => (11,4,0), 58 => (1,0,12), 59 => (8,15,0), 60 => (6,6,0), 61 => (12,5,0), 62 => (12,6,0), 63 => (14,8,0), 64 => (14,9,0), 65 => (14,10,0), 66 => (12,5,0), 67 => (11,12,12), 68 => (14,14,14), 69 => (13,14,14), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (15,14,14), 74 => (7,11,10), 75 => (7,14,1), 76 => (10,10,14), 77 => (9,11,13), 78 => (5,5,9), 79 => (5,5,9), 80 => (5,3,11), 81 => (7,12,1), 82 => (8,14,0), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (8,14,0), 88 => (7,12,0), 89 => (4,0,0), 90 => (8,3,1), 91 => (11,7,5), 92 => (12,8,6), 93 => (12,8,6), 94 => (11,7,5), 95 => (11,7,5), 96 => (13,9,7), 97 => (14,10,7), 98 => (14,10,9), 99 => (14,12,11), 100 => (14,9,7), 101 => (12,7,5), 102 => (0,0,0), 103 => (8,4,1), 104 => (12,8,6), 105 => (15,11,9), 106 => (5,2,0), 107 => (8,3,1), 108 => (10,6,4), 109 => (13,9,7), 110 => (11,6,2), 111 => (5,6,15), 112 => (6,6,15), 113 => (11,11,9), 114 => (10,10,9), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (13,13,14), 119 => (11,11,14), 120 => (8,8,15), 121 => (0,0,9), 122 => (0,0,4), 123 => (0,0,10), 124 => (0,0,10), 125 => (0,1,13), 126 => (6,7,14), 127 => (1,2,14), 128 => (0,1,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			50 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,0,3), 33 => (6,6,14), 34 => (11,11,14), 35 => (13,13,14), 36 => (11,10,14), 37 => (3,3,9), 38 => (4,4,5), 39 => (0,0,3), 40 => (0,0,13), 41 => (6,6,14), 42 => (10,10,14), 43 => (13,13,14), 44 => (7,7,10), 45 => (5,5,9), 46 => (5,6,10), 47 => (8,4,2), 48 => (9,9,11), 49 => (6,9,15), 50 => (10,13,15), 51 => (14,7,0), 52 => (13,10,2), 53 => (10,11,12), 54 => (13,10,2), 55 => (14,10,0), 56 => (14,9,0), 57 => (12,6,0), 58 => (7,1,3), 59 => (8,15,0), 60 => (6,5,0), 61 => (13,6,0), 62 => (6,0,0), 63 => (12,6,0), 64 => (14,7,0), 65 => (14,10,0), 66 => (14,8,0), 67 => (11,3,0), 68 => (11,12,11), 69 => (14,14,14), 70 => (14,14,14), 71 => (14,14,14), 72 => (14,14,14), 73 => (9,11,14), 74 => (8,10,14), 75 => (8,11,2), 76 => (6,0,0), 77 => (9,12,15), 78 => (7,7,11), 79 => (6,7,8), 80 => (7,12,1), 81 => (8,14,0), 82 => (8,14,0), 83 => (8,14,0), 84 => (8,14,0), 85 => (8,14,0), 86 => (8,14,0), 87 => (6,12,0), 88 => (7,1,2), 89 => (2,1,0), 90 => (10,6,4), 91 => (12,8,6), 92 => (11,7,5), 93 => (11,7,5), 94 => (13,9,7), 95 => (13,9,7), 96 => (14,10,8), 97 => (14,10,8), 98 => (14,9,7), 99 => (14,9,7), 100 => (14,10,8), 101 => (12,7,3), 102 => (0,0,11), 103 => (0,0,1), 104 => (8,4,1), 105 => (13,9,7), 106 => (1,0,0), 107 => (12,7,5), 108 => (12,8,6), 109 => (12,8,6), 110 => (10,5,2), 111 => (5,6,15), 112 => (5,5,14), 113 => (15,15,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (12,12,14), 117 => (10,10,14), 118 => (6,6,14), 119 => (0,0,13), 120 => (0,0,3), 121 => (4,4,5), 122 => (3,3,9), 123 => (11,10,14), 124 => (13,13,14), 125 => (11,11,14), 126 => (6,6,14), 127 => (0,0,3), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			51 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,1,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,1,10), 33 => (0,0,8), 34 => (10,10,15), 35 => (14,14,14), 36 => (14,14,14), 37 => (15,15,14), 38 => (15,15,14), 39 => (15,15,15), 40 => (15,15,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (9,9,11), 45 => (5,5,9), 46 => (6,6,11), 47 => (7,4,5), 48 => (12,4,0), 49 => (12,8,2), 50 => (9,10,12), 51 => (11,10,8), 52 => (14,9,0), 53 => (12,10,3), 54 => (14,9,0), 55 => (14,10,0), 56 => (14,9,0), 57 => (14,8,0), 58 => (12,4,0), 59 => (8,13,0), 60 => (6,12,0), 61 => (10,4,0), 62 => (9,3,0), 63 => (10,4,0), 64 => (13,7,0), 65 => (14,8,0), 66 => (14,10,0), 67 => (13,7,0), 68 => (10,6,2), 69 => (11,15,15), 70 => (13,15,15), 71 => (14,15,15), 72 => (14,15,15), 73 => (11,15,15), 74 => (8,9,12), 75 => (11,4,0), 76 => (14,9,0), 77 => (6,1,1), 78 => (4,3,9), 79 => (7,14,1), 80 => (7,15,0), 81 => (7,15,0), 82 => (7,15,0), 83 => (7,15,0), 84 => (7,15,0), 85 => (7,15,0), 86 => (6,12,0), 87 => (5,1,1), 88 => (7,4,1), 89 => (2,1,0), 90 => (13,9,7), 91 => (12,9,7), 92 => (14,11,9), 93 => (14,10,8), 94 => (14,10,8), 95 => (14,10,8), 96 => (14,10,8), 97 => (14,10,8), 98 => (14,10,8), 99 => (14,10,8), 100 => (15,11,8), 101 => (5,3,9), 102 => (1,1,15), 103 => (0,0,13), 104 => (0,0,5), 105 => (9,5,0), 106 => (8,4,2), 107 => (9,5,3), 108 => (15,10,8), 109 => (11,7,5), 110 => (12,8,6), 111 => (6,4,6), 112 => (4,5,14), 113 => (15,15,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (15,15,14), 120 => (15,15,15), 121 => (15,15,14), 122 => (15,15,14), 123 => (14,14,14), 124 => (14,14,14), 125 => (10,10,15), 126 => (0,0,8), 127 => (0,1,10), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			52 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,1,14), 11 => (0,1,14), 12 => (4,5,12), 13 => (0,1,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,1,9), 34 => (0,0,8), 35 => (9,9,15), 36 => (13,13,14), 37 => (14,14,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (15,15,14), 45 => (5,5,10), 46 => (1,2,4), 47 => (8,5,6), 48 => (10,4,0), 49 => (11,6,0), 50 => (15,8,0), 51 => (12,9,4), 52 => (14,8,0), 53 => (14,11,0), 54 => (14,11,0), 55 => (14,11,0), 56 => (14,11,0), 57 => (11,7,0), 58 => (8,3,0), 59 => (6,0,0), 60 => (8,8,0), 61 => (10,0,0), 62 => (12,3,0), 63 => (9,0,0), 64 => (12,3,0), 65 => (13,4,0), 66 => (13,4,0), 67 => (10,1,0), 68 => (8,0,0), 69 => (8,0,0), 70 => (8,0,0), 71 => (7,0,0), 72 => (9,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (12,0,0), 76 => (11,0,0), 77 => (12,0,0), 78 => (12,0,0), 79 => (12,0,0), 80 => (12,0,0), 81 => (12,0,0), 82 => (12,0,0), 83 => (12,0,0), 84 => (12,0,0), 85 => (12,0,0), 86 => (12,0,0), 87 => (10,0,0), 88 => (8,0,0), 89 => (9,0,0), 90 => (8,0,0), 91 => (7,0,0), 92 => (10,1,1), 93 => (13,5,4), 94 => (13,5,4), 95 => (13,5,4), 96 => (13,5,4), 97 => (13,5,4), 98 => (13,5,4), 99 => (11,5,4), 100 => (9,5,4), 101 => (3,0,2), 102 => (0,0,9), 103 => (0,0,14), 104 => (0,0,10), 105 => (0,0,11), 106 => (6,3,0), 107 => (4,1,0), 108 => (15,11,9), 109 => (13,9,7), 110 => (12,8,6), 111 => (6,4,6), 112 => (4,5,14), 113 => (15,15,14), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (14,14,14), 123 => (13,13,14), 124 => (9,9,15), 125 => (0,0,8), 126 => (0,1,9), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			53 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,1,14), 10 => (1,2,12), 11 => (5,7,14), 12 => (10,12,14), 13 => (4,5,12), 14 => (0,1,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,1,9), 35 => (0,0,8), 36 => (9,9,15), 37 => (13,13,14), 38 => (14,14,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,14,14), 43 => (14,14,14), 44 => (14,15,15), 45 => (7,8,13), 46 => (4,0,0), 47 => (4,0,0), 48 => (9,5,0), 49 => (12,2,0), 50 => (11,2,0), 51 => (13,4,0), 52 => (13,4,0), 53 => (12,2,0), 54 => (11,0,0), 55 => (11,0,0), 56 => (11,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (12,0,0), 60 => (12,0,0), 61 => (12,0,0), 62 => (11,0,0), 63 => (12,0,0), 64 => (12,0,0), 65 => (12,0,0), 66 => (12,0,0), 67 => (12,0,0), 68 => (12,0,0), 69 => (12,0,0), 70 => (12,0,0), 71 => (12,0,0), 72 => (12,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (12,0,0), 76 => (12,0,0), 77 => (12,0,0), 78 => (12,0,0), 79 => (12,0,0), 80 => (12,0,0), 81 => (12,0,0), 82 => (12,0,0), 83 => (12,0,0), 84 => (12,0,0), 85 => (12,0,0), 86 => (12,0,0), 87 => (12,0,0), 88 => (12,0,0), 89 => (12,0,0), 90 => (12,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (11,0,0), 94 => (12,0,0), 95 => (12,0,0), 96 => (12,0,0), 97 => (12,0,0), 98 => (12,0,0), 99 => (12,0,0), 100 => (12,0,0), 101 => (12,0,0), 102 => (13,0,0), 103 => (13,0,0), 104 => (13,0,0), 105 => (13,0,0), 106 => (8,0,0), 107 => (8,1,0), 108 => (12,4,3), 109 => (13,5,4), 110 => (11,2,0), 111 => (4,7,15), 112 => (4,5,15), 113 => (15,15,15), 114 => (14,14,14), 115 => (14,14,14), 116 => (14,14,14), 117 => (14,14,14), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (14,14,14), 122 => (13,13,14), 123 => (9,9,15), 124 => (0,0,8), 125 => (0,1,9), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			54 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,1,14), 11 => (0,0,14), 12 => (5,7,14), 13 => (0,1,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,1,9), 36 => (0,0,8), 37 => (10,10,15), 38 => (12,12,14), 39 => (14,14,14), 40 => (14,14,14), 41 => (14,14,14), 42 => (14,15,15), 43 => (14,15,15), 44 => (13,6,6), 45 => (10,3,3), 46 => (12,0,0), 47 => (12,0,0), 48 => (12,0,0), 49 => (12,0,0), 50 => (12,0,0), 51 => (12,0,0), 52 => (12,0,0), 53 => (12,0,0), 54 => (11,0,0), 55 => (12,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (12,0,0), 60 => (11,0,0), 61 => (12,0,0), 62 => (14,9,7), 63 => (14,8,6), 64 => (8,11,15), 65 => (9,10,15), 66 => (9,10,15), 67 => (11,9,11), 68 => (14,8,7), 69 => (13,3,2), 70 => (12,0,0), 71 => (12,0,0), 72 => (12,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (12,0,0), 76 => (7,10,13), 77 => (9,10,15), 78 => (9,10,15), 79 => (9,10,15), 80 => (9,11,15), 81 => (9,0,0), 82 => (12,0,0), 83 => (12,0,0), 84 => (12,0,0), 85 => (10,4,3), 86 => (9,11,15), 87 => (9,10,15), 88 => (9,10,15), 89 => (9,11,15), 90 => (9,4,3), 91 => (12,0,0), 92 => (12,0,0), 93 => (13,0,0), 94 => (5,4,3), 95 => (9,11,15), 96 => (9,10,15), 97 => (9,10,15), 98 => (9,10,15), 99 => (9,11,15), 100 => (9,4,3), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (12,0,0), 107 => (12,0,0), 108 => (11,0,0), 109 => (12,0,0), 110 => (12,0,0), 111 => (13,0,0), 112 => (13,0,0), 113 => (11,0,0), 114 => (13,7,7), 115 => (12,5,5), 116 => (14,15,15), 117 => (14,15,15), 118 => (14,14,14), 119 => (14,14,14), 120 => (14,14,14), 121 => (12,12,14), 122 => (10,10,15), 123 => (0,0,8), 124 => (0,1,9), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			55 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,1,14), 12 => (1,2,12), 13 => (0,1,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,1,9), 37 => (0,0,8), 38 => (5,5,14), 39 => (11,11,14), 40 => (13,14,14), 41 => (14,11,11), 42 => (12,2,2), 43 => (11,0,0), 44 => (11,0,0), 45 => (12,0,0), 46 => (13,4,3), 47 => (14,8,6), 48 => (8,11,15), 49 => (9,10,15), 50 => (9,10,15), 51 => (9,10,15), 52 => (9,10,15), 53 => (11,9,11), 54 => (14,9,7), 55 => (13,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (11,0,0), 60 => (13,3,2), 61 => (9,11,15), 62 => (2,2,14), 63 => (2,3,14), 64 => (3,3,14), 65 => (3,3,14), 66 => (3,3,14), 67 => (2,3,14), 68 => (2,3,14), 69 => (6,7,15), 70 => (11,10,12), 71 => (12,0,0), 72 => (12,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (13,0,0), 76 => (0,1,6), 77 => (4,4,14), 78 => (4,4,14), 79 => (4,4,14), 80 => (4,4,14), 81 => (0,2,7), 82 => (14,0,0), 83 => (12,0,0), 84 => (10,0,0), 85 => (0,0,0), 86 => (5,5,15), 87 => (4,4,14), 88 => (4,4,14), 89 => (4,5,15), 90 => (4,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (5,0,0), 94 => (0,0,0), 95 => (5,5,15), 96 => (4,4,14), 97 => (4,4,14), 98 => (4,4,14), 99 => (4,5,15), 100 => (4,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (12,0,0), 107 => (13,3,2), 108 => (14,8,7), 109 => (11,9,11), 110 => (9,10,15), 111 => (9,10,15), 112 => (8,11,15), 113 => (14,8,6), 114 => (14,7,6), 115 => (14,8,7), 116 => (11,0,0), 117 => (12,2,2), 118 => (14,11,11), 119 => (13,14,14), 120 => (11,11,14), 121 => (5,5,14), 122 => (0,0,8), 123 => (0,1,9), 124 => (0,1,15), 125 => (0,1,14), 126 => (0,1,14), 127 => (0,1,14), 128 => (0,1,14), 129 => (0,2,14), 130 => (0,1,14), 131 => (0,1,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			56 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,1,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,1,10), 38 => (0,0,3), 39 => (5,5,15), 40 => (10,7,11), 41 => (6,0,0), 42 => (12,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (9,0,0), 46 => (0,2,11), 47 => (2,3,15), 48 => (3,3,14), 49 => (3,3,14), 50 => (3,3,14), 51 => (3,3,14), 52 => (3,3,14), 53 => (2,3,14), 54 => (2,4,15), 55 => (1,0,0), 56 => (13,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (13,0,0), 60 => (5,7,11), 61 => (5,5,14), 62 => (6,6,14), 63 => (6,6,14), 64 => (6,6,14), 65 => (6,6,14), 66 => (6,6,14), 67 => (6,6,14), 68 => (6,6,14), 69 => (5,5,14), 70 => (6,7,15), 71 => (7,5,7), 72 => (13,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (13,0,0), 76 => (1,2,7), 77 => (6,6,14), 78 => (5,5,14), 79 => (5,5,14), 80 => (5,5,14), 81 => (6,6,15), 82 => (2,0,2), 83 => (14,0,0), 84 => (0,0,0), 85 => (0,0,0), 86 => (6,6,15), 87 => (5,5,14), 88 => (5,5,14), 89 => (5,6,15), 90 => (5,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (6,0,0), 94 => (0,0,0), 95 => (6,6,15), 96 => (5,5,14), 97 => (5,5,14), 98 => (5,5,14), 99 => (5,6,15), 100 => (5,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (13,0,0), 106 => (12,11,12), 107 => (5,7,15), 108 => (2,3,14), 109 => (2,3,14), 110 => (3,3,14), 111 => (3,3,14), 112 => (3,3,14), 113 => (2,3,14), 114 => (2,3,15), 115 => (0,1,7), 116 => (13,0,0), 117 => (12,0,0), 118 => (6,0,0), 119 => (10,7,11), 120 => (5,5,15), 121 => (0,0,3), 122 => (0,1,10), 123 => (0,1,15), 124 => (9,10,5), 125 => (7,8,6), 126 => (9,10,6), 127 => (3,4,6), 128 => (9,10,6), 129 => (0,0,11), 130 => (4,6,11), 131 => (3,4,5), 132 => (0,1,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			57 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,15), 39 => (0,0,4), 40 => (8,0,2), 41 => (4,0,0), 42 => (12,0,0), 43 => (12,0,0), 44 => (9,0,0), 45 => (2,5,12), 46 => (6,6,14), 47 => (6,6,14), 48 => (6,6,14), 49 => (6,6,14), 50 => (6,6,14), 51 => (6,6,14), 52 => (6,6,14), 53 => (6,6,15), 54 => (5,5,11), 55 => (0,0,0), 56 => (5,0,0), 57 => (12,0,0), 58 => (13,0,0), 59 => (2,1,2), 60 => (7,7,15), 61 => (7,7,14), 62 => (7,7,14), 63 => (7,7,14), 64 => (7,7,14), 65 => (7,7,15), 66 => (8,8,15), 67 => (8,8,15), 68 => (7,7,14), 69 => (6,6,14), 70 => (8,8,14), 71 => (4,5,11), 72 => (0,0,0), 73 => (13,0,0), 74 => (11,0,0), 75 => (12,0,0), 76 => (2,4,7), 77 => (8,8,14), 78 => (8,8,14), 79 => (8,8,14), 80 => (8,8,14), 81 => (8,8,14), 82 => (5,6,11), 83 => (10,0,0), 84 => (0,0,0), 85 => (0,0,0), 86 => (9,9,15), 87 => (8,8,14), 88 => (8,8,14), 89 => (8,9,15), 90 => (5,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (6,0,0), 94 => (0,0,0), 95 => (9,9,15), 96 => (8,8,14), 97 => (8,8,14), 98 => (8,8,14), 99 => (8,9,15), 100 => (5,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (14,0,0), 105 => (2,0,2), 106 => (5,6,15), 107 => (5,5,14), 108 => (6,6,14), 109 => (6,6,14), 110 => (6,6,14), 111 => (6,6,14), 112 => (6,6,14), 113 => (6,6,14), 114 => (6,6,14), 115 => (1,3,7), 116 => (13,0,0), 117 => (12,0,0), 118 => (4,0,0), 119 => (8,0,2), 120 => (0,0,4), 121 => (0,2,15), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,0,5), 125 => (8,9,2), 126 => (0,0,2), 127 => (0,0,7), 128 => (7,7,0), 129 => (9,9,2), 130 => (3,3,1), 131 => (8,8,0), 132 => (0,1,15), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			58 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (10,0,0), 41 => (4,0,0), 42 => (12,0,0), 43 => (12,0,0), 44 => (3,1,2), 45 => (7,7,15), 46 => (7,7,14), 47 => (7,7,14), 48 => (7,7,14), 49 => (8,8,15), 50 => (2,2,6), 51 => (3,3,7), 52 => (3,3,7), 53 => (3,3,7), 54 => (1,1,3), 55 => (0,0,0), 56 => (5,0,0), 57 => (13,0,0), 58 => (8,0,0), 59 => (5,6,11), 60 => (8,8,14), 61 => (7,7,14), 62 => (7,7,14), 63 => (8,8,14), 64 => (6,6,11), 65 => (1,1,2), 66 => (0,0,0), 67 => (0,0,0), 68 => (6,6,11), 69 => (8,8,14), 70 => (7,7,14), 71 => (10,10,15), 72 => (0,0,2), 73 => (6,4,3), 74 => (13,7,7), 75 => (14,7,7), 76 => (2,3,6), 77 => (9,9,14), 78 => (9,9,14), 79 => (9,9,14), 80 => (9,9,14), 81 => (9,9,14), 82 => (9,9,15), 83 => (3,4,7), 84 => (0,0,0), 85 => (0,0,0), 86 => (10,10,15), 87 => (9,9,14), 88 => (9,9,14), 89 => (9,10,15), 90 => (4,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (5,0,0), 94 => (0,0,0), 95 => (10,10,15), 96 => (9,9,14), 97 => (9,9,14), 98 => (9,9,14), 99 => (9,10,15), 100 => (4,0,0), 101 => (12,0,0), 102 => (11,0,0), 103 => (13,0,0), 104 => (0,0,0), 105 => (5,6,11), 106 => (7,7,14), 107 => (7,7,14), 108 => (7,7,14), 109 => (7,7,14), 110 => (7,7,14), 111 => (8,8,15), 112 => (8,8,15), 113 => (8,8,15), 114 => (7,8,15), 115 => (5,0,0), 116 => (12,0,0), 117 => (12,0,0), 118 => (4,0,0), 119 => (10,0,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,1,15), 125 => (9,10,6), 126 => (0,0,6), 127 => (0,1,15), 128 => (9,9,0), 129 => (0,0,11), 130 => (0,1,15), 131 => (9,9,0), 132 => (0,1,15), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			59 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (10,0,0), 41 => (5,0,0), 42 => (12,0,0), 43 => (13,0,0), 44 => (2,4,7), 45 => (8,8,14), 46 => (7,7,14), 47 => (7,7,14), 48 => (8,8,14), 49 => (3,3,5), 50 => (0,0,0), 51 => (0,0,0), 52 => (0,0,0), 53 => (0,0,0), 54 => (0,0,0), 55 => (0,0,0), 56 => (5,2,2), 57 => (14,7,7), 58 => (5,2,1), 59 => (10,11,15), 60 => (10,10,14), 61 => (10,10,14), 62 => (10,10,14), 63 => (9,9,12), 64 => (0,0,0), 65 => (0,0,0), 66 => (7,7,7), 67 => (7,7,7), 68 => (1,1,0), 69 => (11,11,15), 70 => (10,10,14), 71 => (13,13,14), 72 => (4,4,6), 73 => (0,0,0), 74 => (15,15,15), 75 => (15,15,15), 76 => (3,3,5), 77 => (10,10,14), 78 => (10,10,14), 79 => (10,10,14), 80 => (10,10,14), 81 => (10,10,14), 82 => (10,10,14), 83 => (11,11,15), 84 => (1,1,2), 85 => (0,0,0), 86 => (11,11,15), 87 => (10,10,14), 88 => (10,10,14), 89 => (10,10,14), 90 => (5,6,6), 91 => (15,15,15), 92 => (15,15,15), 93 => (7,7,7), 94 => (0,0,0), 95 => (11,11,15), 96 => (10,10,14), 97 => (10,10,14), 98 => (10,10,14), 99 => (10,10,15), 100 => (5,2,1), 101 => (13,7,7), 102 => (13,7,7), 103 => (6,4,3), 104 => (0,0,2), 105 => (8,8,15), 106 => (7,7,14), 107 => (7,7,14), 108 => (7,7,14), 109 => (9,9,15), 110 => (3,3,6), 111 => (0,0,0), 112 => (0,0,0), 113 => (0,0,0), 114 => (3,5,8), 115 => (9,0,0), 116 => (12,0,0), 117 => (12,0,0), 118 => (5,0,0), 119 => (10,0,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,0,10), 126 => (0,1,10), 127 => (0,2,15), 128 => (0,0,5), 129 => (0,2,15), 130 => (0,2,14), 131 => (0,0,5), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			60 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (10,0,0), 41 => (3,0,0), 42 => (13,0,0), 43 => (12,0,0), 44 => (3,5,7), 45 => (10,10,14), 46 => (10,10,14), 47 => (10,10,14), 48 => (10,10,14), 49 => (8,8,11), 50 => (0,0,0), 51 => (3,3,2), 52 => (7,7,6), 53 => (15,15,15), 54 => (15,15,15), 55 => (15,15,15), 56 => (14,15,15), 57 => (15,15,15), 58 => (2,3,5), 59 => (10,10,14), 60 => (10,10,14), 61 => (10,10,14), 62 => (11,11,15), 63 => (0,0,0), 64 => (2,2,2), 65 => (15,15,15), 66 => (14,14,14), 67 => (15,15,15), 68 => (6,6,5), 69 => (10,10,14), 70 => (10,10,14), 71 => (9,9,14), 72 => (14,14,15), 73 => (0,0,0), 74 => (6,6,6), 75 => (15,15,15), 76 => (3,3,5), 77 => (10,10,14), 78 => (9,9,14), 79 => (9,9,14), 80 => (10,10,14), 81 => (9,9,14), 82 => (9,9,14), 83 => (10,10,14), 84 => (8,8,11), 85 => (0,0,0), 86 => (10,10,15), 87 => (9,9,14), 88 => (9,9,14), 89 => (11,11,15), 90 => (5,5,5), 91 => (14,14,14), 92 => (14,14,14), 93 => (7,7,7), 94 => (0,0,0), 95 => (10,10,15), 96 => (9,9,14), 97 => (9,9,14), 98 => (9,9,14), 99 => (9,9,14), 100 => (5,6,5), 101 => (15,15,15), 102 => (15,15,15), 103 => (0,0,0), 104 => (4,4,6), 105 => (10,10,14), 106 => (10,10,14), 107 => (10,10,14), 108 => (11,11,15), 109 => (0,0,0), 110 => (6,7,6), 111 => (15,7,7), 112 => (15,7,7), 113 => (0,0,0), 114 => (0,0,0), 115 => (13,0,0), 116 => (11,0,0), 117 => (13,0,0), 118 => (3,0,0), 119 => (10,0,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			61 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (10,0,0), 41 => (1,0,0), 42 => (5,0,6), 43 => (15,8,7), 44 => (5,1,0), 45 => (12,13,15), 46 => (9,9,14), 47 => (9,9,14), 48 => (9,9,14), 49 => (9,9,14), 50 => (10,10,15), 51 => (10,10,15), 52 => (10,10,15), 53 => (2,2,4), 54 => (3,3,4), 55 => (11,11,10), 56 => (15,15,15), 57 => (14,14,14), 58 => (6,6,5), 59 => (13,13,15), 60 => (9,9,14), 61 => (10,10,15), 62 => (5,5,6), 63 => (0,0,0), 64 => (11,11,11), 65 => (14,14,14), 66 => (14,14,14), 67 => (15,15,15), 68 => (5,5,5), 69 => (11,11,15), 70 => (9,9,14), 71 => (9,9,14), 72 => (15,15,15), 73 => (0,0,0), 74 => (7,7,7), 75 => (15,15,15), 76 => (6,6,6), 77 => (13,13,15), 78 => (12,12,14), 79 => (12,13,15), 80 => (9,9,10), 81 => (15,15,15), 82 => (13,14,15), 83 => (12,12,14), 84 => (13,13,15), 85 => (9,10,11), 86 => (14,14,15), 87 => (15,15,15), 88 => (15,15,15), 89 => (14,13,11), 90 => (5,5,5), 91 => (14,14,14), 92 => (14,14,14), 93 => (7,7,7), 94 => (0,0,0), 95 => (15,15,15), 96 => (12,12,14), 97 => (12,12,14), 98 => (12,12,15), 99 => (15,15,15), 100 => (5,5,5), 101 => (15,15,15), 102 => (6,6,6), 103 => (0,0,0), 104 => (11,11,15), 105 => (10,10,14), 106 => (10,10,14), 107 => (10,10,14), 108 => (3,3,5), 109 => (11,11,10), 110 => (15,15,15), 111 => (14,14,14), 112 => (14,14,14), 113 => (15,15,15), 114 => (15,15,15), 115 => (13,7,6), 116 => (14,8,7), 117 => (5,0,6), 118 => (1,0,0), 119 => (10,0,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			62 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (10,0,0), 41 => (5,0,0), 42 => (0,0,14), 43 => (13,13,15), 44 => (7,8,15), 45 => (0,0,2), 46 => (15,15,15), 47 => (14,14,15), 48 => (12,13,15), 49 => (14,14,15), 50 => (15,15,15), 51 => (13,14,15), 52 => (12,12,14), 53 => (13,13,15), 54 => (15,15,15), 55 => (1,1,1), 56 => (1,1,1), 57 => (15,15,15), 58 => (2,1,0), 59 => (11,9,7), 60 => (15,15,11), 61 => (15,15,12), 62 => (5,4,3), 63 => (0,0,0), 64 => (15,15,15), 65 => (14,14,14), 66 => (15,15,15), 67 => (10,11,11), 68 => (6,4,1), 69 => (15,15,11), 70 => (15,15,15), 71 => (15,15,15), 72 => (14,8,0), 73 => (0,0,0), 74 => (7,7,7), 75 => (15,15,15), 76 => (1,0,0), 77 => (11,7,2), 78 => (10,8,7), 79 => (11,7,2), 80 => (2,0,0), 81 => (1,0,0), 82 => (9,4,0), 83 => (10,8,7), 84 => (10,8,7), 85 => (10,8,8), 86 => (8,4,0), 87 => (4,0,0), 88 => (4,0,0), 89 => (6,1,0), 90 => (6,6,7), 91 => (14,14,14), 92 => (14,14,14), 93 => (7,7,7), 94 => (0,0,0), 95 => (9,4,0), 96 => (10,8,7), 97 => (10,8,7), 98 => (10,7,2), 99 => (5,0,0), 100 => (6,6,7), 101 => (15,15,15), 102 => (7,7,7), 103 => (0,0,0), 104 => (14,14,15), 105 => (9,9,14), 106 => (9,9,14), 107 => (11,11,15), 108 => (0,0,0), 109 => (15,15,15), 110 => (14,14,14), 111 => (14,14,14), 112 => (14,14,14), 113 => (11,11,15), 114 => (0,0,9), 115 => (7,7,14), 116 => (13,13,15), 117 => (0,0,14), 118 => (5,0,0), 119 => (10,0,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			63 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,15), 40 => (15,1,0), 41 => (0,0,0), 42 => (0,0,13), 43 => (0,0,11), 44 => (0,0,11), 45 => (13,13,15), 46 => (0,0,0), 47 => (1,0,0), 48 => (5,2,0), 49 => (3,0,0), 50 => (3,0,0), 51 => (9,4,0), 52 => (10,8,7), 53 => (10,8,7), 54 => (10,6,2), 55 => (6,3,0), 56 => (0,0,0), 57 => (15,15,15), 58 => (6,6,7), 59 => (5,0,0), 60 => (4,0,0), 61 => (4,0,0), 62 => (4,0,0), 63 => (0,0,0), 64 => (15,15,15), 65 => (15,15,15), 66 => (5,6,7), 67 => (2,0,0), 68 => (5,1,0), 69 => (4,0,0), 70 => (4,0,0), 71 => (5,0,0), 72 => (1,0,0), 73 => (0,0,0), 74 => (6,6,6), 75 => (15,15,15), 76 => (2,0,0), 77 => (5,0,0), 78 => (5,0,0), 79 => (5,0,0), 80 => (4,2,0), 81 => (0,0,0), 82 => (6,2,0), 83 => (4,0,0), 84 => (4,0,0), 85 => (6,2,0), 86 => (7,3,0), 87 => (7,3,0), 88 => (7,3,0), 89 => (9,4,0), 90 => (5,6,7), 91 => (14,14,14), 92 => (14,14,14), 93 => (7,7,7), 94 => (0,0,0), 95 => (7,2,0), 96 => (4,0,0), 97 => (5,0,0), 98 => (4,0,0), 99 => (8,3,0), 100 => (6,6,7), 101 => (15,15,15), 102 => (7,7,7), 103 => (0,0,0), 104 => (12,10,7), 105 => (15,15,11), 106 => (15,15,15), 107 => (15,15,15), 108 => (5,6,6), 109 => (14,14,14), 110 => (14,14,14), 111 => (14,14,14), 112 => (15,15,15), 113 => (4,3,1), 114 => (3,3,6), 115 => (0,0,12), 116 => (0,0,11), 117 => (0,0,13), 118 => (0,0,0), 119 => (15,1,0), 120 => (0,2,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			64 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,1,15), 40 => (11,5,0), 41 => (0,0,0), 42 => (0,0,13), 43 => (0,0,12), 44 => (13,13,14), 45 => (15,15,15), 46 => (15,15,15), 47 => (2,2,3), 48 => (0,0,0), 49 => (0,0,0), 50 => (0,0,0), 51 => (7,2,0), 52 => (4,0,0), 53 => (4,0,0), 54 => (7,3,0), 55 => (11,6,0), 56 => (0,0,0), 57 => (6,6,6), 58 => (11,11,12), 59 => (7,3,0), 60 => (7,3,0), 61 => (7,3,0), 62 => (9,5,0), 63 => (8,4,0), 64 => (2,0,0), 65 => (2,0,0), 66 => (10,6,0), 67 => (9,5,0), 68 => (7,3,0), 69 => (7,3,0), 70 => (7,3,0), 71 => (8,4,0), 72 => (2,1,0), 73 => (0,0,0), 74 => (11,11,11), 75 => (15,15,15), 76 => (4,2,0), 77 => (10,6,0), 78 => (10,6,0), 79 => (10,6,0), 80 => (6,4,0), 81 => (0,0,0), 82 => (1,0,0), 83 => (14,9,0), 84 => (9,5,0), 85 => (9,5,0), 86 => (12,8,0), 87 => (12,8,0), 88 => (12,8,0), 89 => (14,9,0), 90 => (5,5,7), 91 => (14,14,14), 92 => (14,14,14), 93 => (7,7,7), 94 => (0,0,0), 95 => (12,8,0), 96 => (9,5,0), 97 => (10,6,0), 98 => (9,5,0), 99 => (13,8,0), 100 => (5,6,7), 101 => (15,15,15), 102 => (6,6,6), 103 => (0,0,0), 104 => (2,0,0), 105 => (4,0,0), 106 => (4,0,0), 107 => (4,0,0), 108 => (2,2,2), 109 => (15,15,15), 110 => (15,15,15), 111 => (10,11,11), 112 => (2,1,2), 113 => (6,0,0), 114 => (4,3,2), 115 => (15,15,15), 116 => (0,0,12), 117 => (0,0,13), 118 => (0,0,0), 119 => (11,5,0), 120 => (0,1,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			65 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,1,15), 40 => (4,3,3), 41 => (0,0,0), 42 => (0,0,13), 43 => (0,0,12), 44 => (15,15,15), 45 => (0,0,0), 46 => (5,3,0), 47 => (6,4,0), 48 => (7,5,0), 49 => (6,4,0), 50 => (11,8,0), 51 => (11,7,0), 52 => (9,5,0), 53 => (9,5,0), 54 => (10,6,0), 55 => (15,11,0), 56 => (0,0,0), 57 => (7,7,7), 58 => (15,15,15), 59 => (4,3,1), 60 => (15,13,4), 61 => (12,7,0), 62 => (12,8,0), 63 => (12,8,0), 64 => (12,8,0), 65 => (12,8,0), 66 => (12,8,0), 67 => (12,8,0), 68 => (12,8,0), 69 => (12,8,0), 70 => (12,8,0), 71 => (13,9,0), 72 => (0,0,0), 73 => (0,0,0), 74 => (15,15,15), 75 => (14,15,15), 76 => (5,3,0), 77 => (15,11,0), 78 => (14,10,0), 79 => (15,11,0), 80 => (7,4,0), 81 => (0,0,0), 82 => (0,0,0), 83 => (12,9,0), 84 => (14,10,0), 85 => (14,10,0), 86 => (14,13,0), 87 => (14,10,0), 88 => (14,10,0), 89 => (15,10,0), 90 => (5,6,7), 91 => (15,15,15), 92 => (15,15,15), 93 => (7,7,7), 94 => (0,0,0), 95 => (15,11,0), 96 => (14,10,0), 97 => (14,10,0), 98 => (14,10,0), 99 => (15,10,0), 100 => (5,5,7), 101 => (15,15,15), 102 => (11,11,11), 103 => (0,0,0), 104 => (2,1,0), 105 => (11,7,0), 106 => (7,3,0), 107 => (7,3,0), 108 => (11,6,0), 109 => (2,0,0), 110 => (2,0,0), 111 => (6,3,0), 112 => (10,6,0), 113 => (7,3,0), 114 => (1,0,0), 115 => (14,15,15), 116 => (0,0,12), 117 => (0,0,13), 118 => (0,0,0), 119 => (4,3,3), 120 => (0,1,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			66 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,1,15), 40 => (12,8,3), 41 => (0,0,0), 42 => (0,0,13), 43 => (0,0,12), 44 => (0,0,10), 45 => (11,8,0), 46 => (15,10,0), 47 => (14,10,0), 48 => (14,10,0), 49 => (14,10,0), 50 => (14,10,0), 51 => (14,10,0), 52 => (14,10,0), 53 => (14,10,0), 54 => (15,10,0), 55 => (7,6,5), 56 => (0,0,0), 57 => (6,7,7), 58 => (15,15,15), 59 => (15,15,15), 60 => (0,0,2), 61 => (15,15,10), 62 => (15,10,0), 63 => (15,10,0), 64 => (14,10,0), 65 => (14,10,0), 66 => (14,10,0), 67 => (14,10,0), 68 => (15,10,0), 69 => (15,12,3), 70 => (12,11,10), 71 => (0,0,0), 72 => (0,0,0), 73 => (6,4,4), 74 => (13,7,7), 75 => (14,10,7), 76 => (5,7,9), 77 => (15,10,0), 78 => (14,10,0), 79 => (15,10,0), 80 => (7,8,10), 81 => (0,0,0), 82 => (0,0,0), 83 => (0,0,0), 84 => (15,14,10), 85 => (14,13,0), 86 => (14,9,0), 87 => (14,10,0), 88 => (14,10,0), 89 => (15,14,9), 90 => (4,2,2), 91 => (13,7,7), 92 => (13,7,7), 93 => (6,3,3), 94 => (0,0,0), 95 => (15,14,9), 96 => (14,10,0), 97 => (14,10,0), 98 => (14,10,0), 99 => (15,13,8), 100 => (5,6,7), 101 => (15,15,15), 102 => (15,15,15), 103 => (0,0,0), 104 => (0,0,0), 105 => (12,10,5), 106 => (14,9,0), 107 => (12,8,0), 108 => (12,8,0), 109 => (12,8,0), 110 => (12,8,0), 111 => (12,8,0), 112 => (13,9,0), 113 => (15,11,0), 114 => (11,7,0), 115 => (2,2,10), 116 => (0,0,12), 117 => (0,0,13), 118 => (0,0,0), 119 => (12,8,3), 120 => (0,1,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			67 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,1,15), 40 => (15,9,0), 41 => (0,0,2), 42 => (8,8,15), 43 => (6,6,13), 44 => (0,0,5), 45 => (15,15,9), 46 => (15,12,3), 47 => (14,10,0), 48 => (14,10,0), 49 => (14,10,0), 50 => (14,10,0), 51 => (14,10,0), 52 => (14,10,0), 53 => (15,14,9), 54 => (12,11,9), 55 => (0,0,0), 56 => (0,0,0), 57 => (14,0,0), 58 => (11,0,0), 59 => (12,0,0), 60 => (10,0,0), 61 => (0,0,0), 62 => (7,8,9), 63 => (6,6,8), 64 => (15,14,8), 65 => (15,13,8), 66 => (15,14,8), 67 => (11,10,8), 68 => (7,7,9), 69 => (2,3,3), 70 => (0,0,0), 71 => (0,0,0), 72 => (1,0,0), 73 => (13,0,0), 74 => (11,0,0), 75 => (14,5,0), 76 => (0,2,3), 77 => (7,7,9), 78 => (7,7,8), 79 => (7,7,9), 80 => (3,3,3), 81 => (0,0,0), 82 => (12,0,0), 83 => (0,0,0), 84 => (2,2,3), 85 => (7,7,9), 86 => (7,7,8), 87 => (7,7,8), 88 => (7,7,8), 89 => (6,8,8), 90 => (4,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (5,0,0), 94 => (0,0,0), 95 => (7,8,8), 96 => (7,7,8), 97 => (7,7,8), 98 => (7,7,8), 99 => (6,8,8), 100 => (4,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (6,0,0), 104 => (0,0,0), 105 => (0,0,0), 106 => (12,11,10), 107 => (15,12,3), 108 => (15,10,0), 109 => (14,10,0), 110 => (14,10,0), 111 => (14,10,0), 112 => (14,9,0), 113 => (14,10,0), 114 => (15,14,8), 115 => (0,0,5), 116 => (6,6,13), 117 => (8,8,15), 118 => (0,0,2), 119 => (15,9,0), 120 => (0,1,15), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			68 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,15), 39 => (6,0,7), 40 => (14,9,0), 41 => (0,0,0), 42 => (15,15,15), 43 => (15,15,15), 44 => (14,7,7), 45 => (0,0,0), 46 => (1,3,3), 47 => (7,7,9), 48 => (7,7,8), 49 => (7,7,8), 50 => (7,7,8), 51 => (7,7,8), 52 => (7,8,9), 53 => (0,0,0), 54 => (0,0,0), 55 => (1,0,0), 56 => (10,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (12,0,0), 60 => (12,0,0), 61 => (10,0,0), 62 => (1,0,0), 63 => (0,0,0), 64 => (0,0,0), 65 => (0,0,0), 66 => (0,0,0), 67 => (0,0,0), 68 => (0,0,0), 69 => (0,0,0), 70 => (1,0,0), 71 => (10,0,0), 72 => (13,0,0), 73 => (12,0,0), 74 => (12,0,0), 75 => (12,0,0), 76 => (11,6,0), 77 => (0,0,0), 78 => (0,0,0), 79 => (0,0,0), 80 => (0,0,0), 81 => (0,0,0), 82 => (15,0,0), 83 => (1,0,0), 84 => (0,0,0), 85 => (0,0,0), 86 => (0,0,0), 87 => (0,0,0), 88 => (0,0,0), 89 => (0,0,0), 90 => (13,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (5,0,0), 94 => (0,0,0), 95 => (0,0,0), 96 => (0,0,0), 97 => (0,0,0), 98 => (0,0,0), 99 => (0,0,0), 100 => (13,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (13,0,0), 104 => (1,0,0), 105 => (0,0,0), 106 => (0,0,0), 107 => (2,3,3), 108 => (7,7,9), 109 => (11,10,8), 110 => (15,14,8), 111 => (15,13,8), 112 => (15,14,8), 113 => (5,6,8), 114 => (5,7,8), 115 => (10,2,1), 116 => (15,15,15), 117 => (15,15,15), 118 => (0,0,0), 119 => (14,9,0), 120 => (6,0,7), 121 => (0,2,15), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			69 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,15), 36 => (2,1,11), 37 => (6,1,7), 38 => (11,0,0), 39 => (4,0,0), 40 => (14,10,0), 41 => (0,0,0), 42 => (14,3,3), 43 => (11,0,0), 44 => (12,0,0), 45 => (13,0,0), 46 => (5,0,0), 47 => (1,0,0), 48 => (0,0,0), 49 => (0,0,0), 50 => (0,0,0), 51 => (0,0,0), 52 => (0,0,0), 53 => (2,0,0), 54 => (5,0,0), 55 => (13,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (12,0,0), 60 => (11,0,0), 61 => (12,0,0), 62 => (12,0,0), 63 => (14,0,0), 64 => (5,0,0), 65 => (6,0,0), 66 => (6,0,0), 67 => (5,0,0), 68 => (5,0,0), 69 => (15,0,0), 70 => (13,0,0), 71 => (12,0,0), 72 => (12,0,0), 73 => (11,0,0), 74 => (13,0,0), 75 => (11,0,0), 76 => (14,6,0), 77 => (13,0,0), 78 => (14,0,0), 79 => (14,0,0), 80 => (13,0,0), 81 => (13,0,0), 82 => (12,1,0), 83 => (12,5,0), 84 => (12,8,0), 85 => (14,0,0), 86 => (14,0,0), 87 => (13,0,0), 88 => (14,0,0), 89 => (13,0,0), 90 => (12,0,0), 91 => (12,0,0), 92 => (12,0,0), 93 => (12,0,0), 94 => (14,0,0), 95 => (13,0,0), 96 => (14,0,0), 97 => (13,0,0), 98 => (14,0,0), 99 => (14,0,0), 100 => (12,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (13,0,0), 105 => (10,0,0), 106 => (1,0,0), 107 => (0,0,0), 108 => (0,0,0), 109 => (0,0,0), 110 => (0,0,0), 111 => (0,0,0), 112 => (0,0,0), 113 => (1,0,0), 114 => (9,0,0), 115 => (12,0,0), 116 => (11,0,0), 117 => (14,3,3), 118 => (0,0,0), 119 => (14,10,0), 120 => (4,0,0), 121 => (11,0,0), 122 => (6,1,7), 123 => (2,1,11), 124 => (0,2,15), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			70 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,15), 33 => (2,1,11), 34 => (5,1,7), 35 => (14,0,0), 36 => (13,0,0), 37 => (9,0,0), 38 => (5,0,0), 39 => (5,0,0), 40 => (14,10,0), 41 => (0,0,0), 42 => (13,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (12,0,0), 46 => (12,0,0), 47 => (13,0,0), 48 => (13,0,0), 49 => (13,0,0), 50 => (13,0,0), 51 => (13,0,0), 52 => (13,0,0), 53 => (13,0,0), 54 => (12,0,0), 55 => (12,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (11,0,0), 60 => (15,15,15), 61 => (14,15,15), 62 => (15,15,15), 63 => (5,7,7), 64 => (6,7,7), 65 => (6,7,7), 66 => (6,7,7), 67 => (15,15,15), 68 => (6,7,7), 69 => (0,4,4), 70 => (13,0,0), 71 => (12,0,0), 72 => (3,0,0), 73 => (15,15,15), 74 => (0,0,0), 75 => (15,15,15), 76 => (4,5,6), 77 => (11,12,12), 78 => (6,7,7), 79 => (5,7,7), 80 => (11,12,12), 81 => (11,13,13), 82 => (0,1,1), 83 => (11,12,12), 84 => (6,7,7), 85 => (5,7,7), 86 => (5,7,7), 87 => (11,12,12), 88 => (6,7,7), 89 => (6,7,7), 90 => (5,7,7), 91 => (5,7,7), 92 => (5,7,7), 93 => (10,12,12), 94 => (6,7,7), 95 => (11,12,12), 96 => (0,1,1), 97 => (12,13,13), 98 => (5,7,7), 99 => (0,3,3), 100 => (13,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (13,0,0), 107 => (14,0,0), 108 => (5,0,0), 109 => (6,0,0), 110 => (6,0,0), 111 => (5,0,0), 112 => (14,0,0), 113 => (13,0,0), 114 => (12,0,0), 115 => (12,0,0), 116 => (12,0,0), 117 => (13,0,0), 118 => (0,0,0), 119 => (14,10,0), 120 => (5,0,0), 121 => (5,0,0), 122 => (9,0,0), 123 => (13,0,0), 124 => (14,0,0), 125 => (5,1,7), 126 => (2,1,11), 127 => (0,2,15), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			71 => (0 => (0,1,14), 1 => (0,1,14), 2 => (0,1,14), 3 => (0,1,14), 4 => (0,1,14), 5 => (0,1,14), 6 => (0,1,14), 7 => (0,1,14), 8 => (0,1,14), 9 => (0,1,14), 10 => (0,1,14), 11 => (0,1,14), 12 => (0,1,14), 13 => (0,1,14), 14 => (0,1,14), 15 => (0,1,14), 16 => (0,1,14), 17 => (0,1,14), 18 => (0,1,14), 19 => (0,1,14), 20 => (0,1,14), 21 => (0,1,14), 22 => (0,1,14), 23 => (0,1,14), 24 => (0,1,14), 25 => (0,1,14), 26 => (0,1,14), 27 => (0,2,14), 28 => (0,2,15), 29 => (0,2,15), 30 => (2,1,11), 31 => (5,1,7), 32 => (14,0,0), 33 => (13,0,0), 34 => (12,0,0), 35 => (12,0,0), 36 => (12,0,0), 37 => (9,0,0), 38 => (5,0,0), 39 => (5,0,0), 40 => (10,2,0), 41 => (5,0,0), 42 => (12,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (12,0,0), 46 => (12,0,0), 47 => (12,0,0), 48 => (12,0,0), 49 => (12,0,0), 50 => (12,0,0), 51 => (12,0,0), 52 => (12,0,0), 53 => (12,0,0), 54 => (12,0,0), 55 => (12,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (13,0,0), 60 => (0,0,0), 61 => (15,15,15), 62 => (0,0,0), 63 => (6,7,7), 64 => (15,15,15), 65 => (15,15,15), 66 => (5,5,5), 67 => (15,15,15), 68 => (5,6,6), 69 => (5,0,0), 70 => (12,0,0), 71 => (12,0,0), 72 => (4,0,0), 73 => (15,15,15), 74 => (15,15,15), 75 => (14,14,14), 76 => (5,5,5), 77 => (11,11,11), 78 => (0,0,0), 79 => (7,7,7), 80 => (5,5,5), 81 => (5,5,5), 82 => (7,7,7), 83 => (15,15,15), 84 => (0,0,0), 85 => (15,15,15), 86 => (5,5,5), 87 => (11,11,11), 88 => (1,1,1), 89 => (6,6,6), 90 => (15,15,15), 91 => (15,15,15), 92 => (5,5,5), 93 => (15,15,15), 94 => (0,0,0), 95 => (15,15,15), 96 => (7,7,7), 97 => (5,5,5), 98 => (11,11,11), 99 => (6,7,7), 100 => (12,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (12,0,0), 107 => (12,0,0), 108 => (12,0,0), 109 => (12,0,0), 110 => (12,0,0), 111 => (12,0,0), 112 => (12,0,0), 113 => (12,0,0), 114 => (12,0,0), 115 => (12,0,0), 116 => (12,0,0), 117 => (12,0,0), 118 => (5,0,0), 119 => (10,2,0), 120 => (5,0,0), 121 => (5,0,0), 122 => (9,0,0), 123 => (12,0,0), 124 => (12,0,0), 125 => (12,0,0), 126 => (13,0,0), 127 => (14,0,0), 128 => (5,1,7), 129 => (2,1,11), 130 => (0,2,15), 131 => (0,2,15), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,1,14), 135 => (0,1,14), 136 => (0,1,14), 137 => (0,1,14), 138 => (0,1,14), 139 => (0,1,14), 140 => (0,1,14), 141 => (0,1,14), 142 => (0,1,14), 143 => (0,1,14), 144 => (0,1,14), 145 => (0,1,14), 146 => (0,1,14), 147 => (0,1,14), 148 => (0,1,14), 149 => (0,1,14), 150 => (0,1,14), 151 => (0,1,14), 152 => (0,1,14), 153 => (0,1,14), 154 => (0,1,14), 155 => (0,1,14), 156 => (0,1,14), 157 => (0,1,14), 158 => (0,1,14), 159 => (0,1,14)), 
			72 => (0 => (1,3,14), 1 => (1,3,14), 2 => (1,3,14), 3 => (1,3,14), 4 => (1,3,14), 5 => (1,3,14), 6 => (1,3,14), 7 => (1,3,14), 8 => (1,3,14), 9 => (1,3,14), 10 => (1,3,14), 11 => (1,3,14), 12 => (1,3,14), 13 => (1,3,14), 14 => (1,3,14), 15 => (1,3,14), 16 => (1,3,14), 17 => (1,3,14), 18 => (1,3,14), 19 => (1,3,14), 20 => (1,3,14), 21 => (1,3,14), 22 => (1,3,14), 23 => (1,3,14), 24 => (1,3,14), 25 => (0,3,15), 26 => (3,2,11), 27 => (6,1,7), 28 => (9,0,2), 29 => (13,0,0), 30 => (13,0,0), 31 => (12,0,0), 32 => (12,0,0), 33 => (12,0,0), 34 => (12,0,0), 35 => (12,0,0), 36 => (12,0,0), 37 => (9,0,0), 38 => (5,0,0), 39 => (5,0,0), 40 => (9,0,0), 41 => (4,0,0), 42 => (12,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (12,0,0), 46 => (12,0,0), 47 => (12,0,0), 48 => (12,0,0), 49 => (12,0,0), 50 => (12,0,0), 51 => (12,0,0), 52 => (12,0,0), 53 => (12,0,0), 54 => (12,0,0), 55 => (12,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (12,0,0), 60 => (4,0,0), 61 => (15,15,15), 62 => (4,0,0), 63 => (7,8,8), 64 => (6,7,7), 65 => (6,7,7), 66 => (6,7,7), 67 => (15,15,15), 68 => (15,15,15), 69 => (5,8,8), 70 => (12,0,0), 71 => (12,0,0), 72 => (3,0,0), 73 => (15,15,15), 74 => (0,0,0), 75 => (15,15,15), 76 => (5,6,6), 77 => (15,15,15), 78 => (15,15,15), 79 => (5,6,6), 80 => (15,15,15), 81 => (15,15,15), 82 => (0,0,1), 83 => (11,11,11), 84 => (15,15,15), 85 => (15,15,15), 86 => (5,6,6), 87 => (11,12,12), 88 => (7,7,7), 89 => (7,7,7), 90 => (6,7,7), 91 => (6,7,7), 92 => (6,7,7), 93 => (10,11,11), 94 => (15,15,15), 95 => (11,11,11), 96 => (0,1,1), 97 => (15,15,15), 98 => (15,15,15), 99 => (5,7,7), 100 => (12,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (12,0,0), 107 => (12,0,0), 108 => (12,0,0), 109 => (12,0,0), 110 => (12,0,0), 111 => (12,0,0), 112 => (12,0,0), 113 => (12,0,0), 114 => (12,0,0), 115 => (12,0,0), 116 => (12,0,0), 117 => (12,0,0), 118 => (4,0,0), 119 => (9,0,0), 120 => (5,0,0), 121 => (5,0,0), 122 => (9,0,0), 123 => (12,0,0), 124 => (12,0,0), 125 => (12,0,0), 126 => (12,0,0), 127 => (12,0,0), 128 => (12,0,0), 129 => (13,0,0), 130 => (13,0,0), 131 => (10,1,2), 132 => (6,1,7), 133 => (2,2,11), 134 => (0,3,15), 135 => (1,3,14), 136 => (1,3,14), 137 => (1,3,14), 138 => (1,3,14), 139 => (1,3,14), 140 => (1,3,14), 141 => (1,3,14), 142 => (1,3,14), 143 => (1,3,14), 144 => (1,3,14), 145 => (1,3,14), 146 => (1,3,14), 147 => (1,3,14), 148 => (1,3,14), 149 => (1,3,14), 150 => (1,3,14), 151 => (1,3,14), 152 => (1,3,14), 153 => (1,3,14), 154 => (1,3,14), 155 => (1,3,14), 156 => (1,3,14), 157 => (1,3,14), 158 => (1,3,14), 159 => (1,3,14)), 
			73 => (0 => (1,3,14), 1 => (1,3,14), 2 => (1,3,14), 3 => (1,3,14), 4 => (1,3,14), 5 => (1,3,14), 6 => (1,3,14), 7 => (1,3,14), 8 => (1,3,14), 9 => (1,3,14), 10 => (1,3,14), 11 => (1,3,14), 12 => (1,3,14), 13 => (1,3,14), 14 => (1,3,14), 15 => (1,3,14), 16 => (1,3,14), 17 => (1,3,14), 18 => (1,3,14), 19 => (1,3,14), 20 => (1,3,14), 21 => (1,3,14), 22 => (1,3,14), 23 => (1,3,14), 24 => (0,3,15), 25 => (12,0,0), 26 => (13,0,0), 27 => (12,0,0), 28 => (12,0,0), 29 => (12,0,0), 30 => (12,0,0), 31 => (12,0,0), 32 => (12,0,0), 33 => (12,0,0), 34 => (12,0,0), 35 => (11,0,0), 36 => (12,0,0), 37 => (8,0,0), 38 => (7,1,0), 39 => (12,8,0), 40 => (10,1,0), 41 => (4,0,0), 42 => (10,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (12,0,0), 46 => (12,0,0), 47 => (12,0,0), 48 => (12,0,0), 49 => (12,0,0), 50 => (12,0,0), 51 => (12,0,0), 52 => (12,0,0), 53 => (12,0,0), 54 => (12,0,0), 55 => (12,0,0), 56 => (12,0,0), 57 => (12,0,0), 58 => (12,0,0), 59 => (13,0,0), 60 => (10,0,0), 61 => (4,0,0), 62 => (10,0,0), 63 => (5,0,0), 64 => (5,0,0), 65 => (5,0,0), 66 => (5,0,0), 67 => (4,0,0), 68 => (4,0,0), 69 => (4,0,0), 70 => (13,0,0), 71 => (12,0,0), 72 => (9,0,0), 73 => (4,0,0), 74 => (6,0,0), 75 => (4,0,0), 76 => (5,0,0), 77 => (4,0,0), 78 => (3,0,0), 79 => (5,0,0), 80 => (3,0,0), 81 => (3,2,0), 82 => (12,9,0), 83 => (3,0,0), 84 => (4,0,0), 85 => (4,0,0), 86 => (5,0,0), 87 => (5,0,0), 88 => (5,0,0), 89 => (5,0,0), 90 => (5,0,0), 91 => (5,0,0), 92 => (5,0,0), 93 => (5,0,0), 94 => (4,0,0), 95 => (5,0,0), 96 => (10,0,0), 97 => (4,0,0), 98 => (4,0,0), 99 => (5,0,0), 100 => (13,0,0), 101 => (12,0,0), 102 => (12,0,0), 103 => (12,0,0), 104 => (12,0,0), 105 => (12,0,0), 106 => (12,0,0), 107 => (12,0,0), 108 => (12,0,0), 109 => (12,0,0), 110 => (12,0,0), 111 => (12,0,0), 112 => (12,0,0), 113 => (12,0,0), 114 => (12,0,0), 115 => (12,0,0), 116 => (12,0,0), 117 => (10,0,0), 118 => (4,0,0), 119 => (10,1,0), 120 => (12,8,0), 121 => (7,1,0), 122 => (8,0,0), 123 => (12,0,0), 124 => (11,0,0), 125 => (12,0,0), 126 => (12,0,0), 127 => (12,0,0), 128 => (12,0,0), 129 => (12,0,0), 130 => (12,0,0), 131 => (12,0,0), 132 => (12,0,0), 133 => (13,0,0), 134 => (11,0,0), 135 => (0,3,15), 136 => (1,3,14), 137 => (1,3,14), 138 => (1,3,14), 139 => (1,3,14), 140 => (1,3,14), 141 => (1,3,14), 142 => (1,3,14), 143 => (1,3,14), 144 => (1,3,14), 145 => (1,3,14), 146 => (1,3,14), 147 => (1,3,14), 148 => (1,3,14), 149 => (1,3,14), 150 => (1,3,14), 151 => (1,3,14), 152 => (1,3,14), 153 => (1,3,14), 154 => (1,3,14), 155 => (1,3,14), 156 => (1,3,14), 157 => (1,3,14), 158 => (1,3,14), 159 => (1,3,14)), 
			74 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,3,15), 26 => (10,0,1), 27 => (12,0,0), 28 => (12,0,0), 29 => (12,0,0), 30 => (12,0,0), 31 => (12,0,0), 32 => (11,0,0), 33 => (11,0,0), 34 => (11,0,0), 35 => (13,7,7), 36 => (13,11,12), 37 => (14,13,8), 38 => (15,10,0), 39 => (12,8,0), 40 => (11,2,0), 41 => (5,0,0), 42 => (8,0,0), 43 => (12,0,0), 44 => (12,0,0), 45 => (12,0,0), 46 => (12,0,0), 47 => (12,0,0), 48 => (13,0,0), 49 => (13,0,0), 50 => (13,0,0), 51 => (13,0,0), 52 => (5,1,7), 53 => (6,1,7), 54 => (6,1,7), 55 => (6,1,7), 56 => (6,1,7), 57 => (6,1,7), 58 => (8,1,1), 59 => (5,3,12), 60 => (1,2,15), 61 => (8,6,7), 62 => (5,1,0), 63 => (5,1,0), 64 => (5,1,0), 65 => (8,4,0), 66 => (7,4,0), 67 => (7,4,0), 68 => (7,4,0), 69 => (7,4,0), 70 => (7,4,0), 71 => (7,4,0), 72 => (7,4,0), 73 => (7,4,0), 74 => (7,4,0), 75 => (7,4,0), 76 => (7,4,0), 77 => (7,3,0), 78 => (8,4,0), 79 => (13,8,0), 80 => (13,4,0), 81 => (13,4,0), 82 => (13,3,0), 83 => (7,3,0), 84 => (7,4,0), 85 => (7,4,0), 86 => (7,4,0), 87 => (7,4,0), 88 => (7,4,0), 89 => (7,4,0), 90 => (7,4,0), 91 => (7,4,0), 92 => (7,4,0), 93 => (7,4,0), 94 => (8,4,0), 95 => (5,1,0), 96 => (5,1,0), 97 => (5,1,0), 98 => (8,6,7), 99 => (1,2,15), 100 => (5,3,12), 101 => (8,1,1), 102 => (6,1,7), 103 => (6,1,7), 104 => (6,1,7), 105 => (6,1,7), 106 => (6,1,7), 107 => (5,1,7), 108 => (13,0,0), 109 => (13,0,0), 110 => (13,0,0), 111 => (13,0,0), 112 => (12,0,0), 113 => (12,0,0), 114 => (12,0,0), 115 => (12,0,0), 116 => (12,0,0), 117 => (8,0,0), 118 => (5,0,0), 119 => (11,2,0), 120 => (12,8,0), 121 => (15,10,0), 122 => (14,13,8), 123 => (13,11,12), 124 => (13,7,7), 125 => (11,0,0), 126 => (11,0,0), 127 => (11,0,0), 128 => (12,0,0), 129 => (12,0,0), 130 => (12,0,0), 131 => (12,0,0), 132 => (12,0,0), 133 => (10,0,1), 134 => (0,3,15), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			75 => (0 => (2,4,14), 1 => (2,4,14), 2 => (2,4,14), 3 => (2,4,14), 4 => (2,4,14), 5 => (2,4,14), 6 => (2,4,14), 7 => (2,4,14), 8 => (2,4,14), 9 => (2,4,14), 10 => (2,4,14), 11 => (2,4,14), 12 => (2,4,14), 13 => (2,4,14), 14 => (2,4,14), 15 => (2,4,14), 16 => (2,4,14), 17 => (2,4,14), 18 => (2,4,14), 19 => (2,4,14), 20 => (2,4,14), 21 => (2,4,14), 22 => (2,4,14), 23 => (2,4,14), 24 => (2,4,14), 25 => (2,4,14), 26 => (0,4,15), 27 => (10,0,1), 28 => (12,0,0), 29 => (11,0,0), 30 => (11,0,0), 31 => (11,0,0), 32 => (13,7,7), 33 => (13,11,11), 34 => (14,15,15), 35 => (14,14,14), 36 => (14,14,15), 37 => (14,12,7), 38 => (14,10,0), 39 => (11,8,0), 40 => (11,2,0), 41 => (4,0,0), 42 => (9,0,0), 43 => (13,0,0), 44 => (13,0,0), 45 => (7,0,0), 46 => (11,0,0), 47 => (3,3,12), 48 => (0,4,15), 49 => (0,4,15), 50 => (0,4,15), 51 => (0,4,15), 52 => (1,4,14), 53 => (1,4,14), 54 => (1,4,14), 55 => (1,4,14), 56 => (1,4,14), 57 => (1,4,15), 58 => (0,2,10), 59 => (2,2,4), 60 => (5,5,15), 61 => (0,0,13), 62 => (5,5,11), 63 => (10,7,2), 64 => (13,8,0), 65 => (12,7,0), 66 => (12,7,0), 67 => (12,7,0), 68 => (12,7,0), 69 => (12,7,0), 70 => (12,7,0), 71 => (12,7,0), 72 => (12,7,0), 73 => (12,8,0), 74 => (13,8,0), 75 => (13,8,0), 76 => (13,8,0), 77 => (12,8,0), 78 => (15,15,0), 79 => (15,15,3), 80 => (15,15,8), 81 => (15,15,3), 82 => (15,15,0), 83 => (14,9,0), 84 => (13,8,0), 85 => (13,8,0), 86 => (12,8,0), 87 => (12,7,0), 88 => (12,7,0), 89 => (12,7,0), 90 => (12,7,0), 91 => (12,7,0), 92 => (12,7,0), 93 => (12,7,0), 94 => (12,7,0), 95 => (13,8,0), 96 => (10,7,2), 97 => (5,5,11), 98 => (0,0,13), 99 => (5,5,15), 100 => (2,2,4), 101 => (0,2,10), 102 => (1,4,15), 103 => (1,4,14), 104 => (1,4,14), 105 => (1,4,14), 106 => (1,4,14), 107 => (1,4,14), 108 => (0,4,15), 109 => (0,4,15), 110 => (0,4,15), 111 => (0,4,15), 112 => (3,3,12), 113 => (11,0,0), 114 => (7,0,0), 115 => (13,0,0), 116 => (13,0,0), 117 => (9,0,0), 118 => (4,0,0), 119 => (11,2,0), 120 => (11,8,0), 121 => (14,10,0), 122 => (14,12,7), 123 => (14,14,15), 124 => (14,14,14), 125 => (14,15,15), 126 => (13,11,11), 127 => (13,7,7), 128 => (11,0,0), 129 => (11,0,0), 130 => (11,0,0), 131 => (12,0,0), 132 => (10,0,1), 133 => (0,4,15), 134 => (2,4,14), 135 => (2,4,14), 136 => (2,4,14), 137 => (2,4,14), 138 => (2,4,14), 139 => (2,4,14), 140 => (2,4,14), 141 => (2,4,14), 142 => (2,4,14), 143 => (2,4,14), 144 => (2,4,14), 145 => (2,4,14), 146 => (2,4,14), 147 => (2,4,14), 148 => (2,4,14), 149 => (2,4,14), 150 => (2,4,14), 151 => (2,4,14), 152 => (2,4,14), 153 => (2,4,14), 154 => (2,4,14), 155 => (2,4,14), 156 => (2,4,14), 157 => (2,4,14), 158 => (2,4,14), 159 => (2,4,14)), 
			76 => (0 => (2,4,14), 1 => (2,4,14), 2 => (2,4,14), 3 => (2,4,14), 4 => (2,4,14), 5 => (2,4,14), 6 => (2,4,14), 7 => (2,4,14), 8 => (2,4,14), 9 => (2,4,14), 10 => (2,4,14), 11 => (2,4,14), 12 => (2,4,14), 13 => (2,4,14), 14 => (2,4,14), 15 => (2,4,14), 16 => (2,4,14), 17 => (2,4,14), 18 => (2,4,14), 19 => (2,4,14), 20 => (2,4,14), 21 => (2,4,14), 22 => (2,4,14), 23 => (2,4,14), 24 => (2,4,14), 25 => (2,4,14), 26 => (2,4,14), 27 => (0,4,15), 28 => (10,0,0), 29 => (13,8,7), 30 => (13,11,11), 31 => (14,15,15), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,12,7), 38 => (14,10,0), 39 => (11,8,0), 40 => (10,4,0), 41 => (7,0,0), 42 => (6,0,0), 43 => (0,0,0), 44 => (0,0,0), 45 => (3,1,0), 46 => (10,0,0), 47 => (0,4,15), 48 => (2,4,14), 49 => (2,4,14), 50 => (2,4,14), 51 => (2,4,14), 52 => (2,4,14), 53 => (2,4,14), 54 => (2,4,14), 55 => (2,4,14), 56 => (2,4,14), 57 => (2,4,14), 58 => (2,4,14), 59 => (1,4,15), 60 => (1,1,3), 61 => (6,6,15), 62 => (2,2,14), 63 => (0,1,14), 64 => (12,10,7), 65 => (15,15,0), 66 => (14,15,0), 67 => (14,14,0), 68 => (14,14,0), 69 => (14,14,0), 70 => (14,14,0), 71 => (14,14,0), 72 => (15,15,3), 73 => (11,11,7), 74 => (5,6,7), 75 => (6,6,7), 76 => (6,6,7), 77 => (5,6,7), 78 => (5,5,7), 79 => (5,5,6), 80 => (5,5,6), 81 => (5,5,6), 82 => (5,5,7), 83 => (5,6,7), 84 => (6,6,7), 85 => (6,6,7), 86 => (11,11,7), 87 => (15,15,3), 88 => (14,14,0), 89 => (14,14,0), 90 => (14,14,0), 91 => (14,14,0), 92 => (14,14,0), 93 => (14,15,0), 94 => (15,15,0), 95 => (12,10,7), 96 => (0,1,14), 97 => (2,2,14), 98 => (6,6,15), 99 => (1,1,3), 100 => (1,4,15), 101 => (2,4,14), 102 => (2,4,14), 103 => (2,4,14), 104 => (2,4,14), 105 => (2,4,14), 106 => (2,4,14), 107 => (2,4,14), 108 => (2,4,14), 109 => (2,4,14), 110 => (2,4,14), 111 => (2,4,14), 112 => (0,4,15), 113 => (10,0,0), 114 => (3,1,0), 115 => (0,0,0), 116 => (0,0,0), 117 => (6,0,0), 118 => (7,0,0), 119 => (10,4,0), 120 => (11,8,0), 121 => (14,10,0), 122 => (14,12,7), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,15,15), 129 => (13,11,11), 130 => (13,8,7), 131 => (10,0,0), 132 => (0,4,15), 133 => (2,4,14), 134 => (2,4,14), 135 => (2,4,14), 136 => (2,4,14), 137 => (2,4,14), 138 => (2,4,14), 139 => (2,4,14), 140 => (2,4,14), 141 => (2,4,14), 142 => (2,4,14), 143 => (2,4,14), 144 => (2,4,14), 145 => (2,4,14), 146 => (2,4,14), 147 => (2,4,14), 148 => (2,4,14), 149 => (2,4,14), 150 => (2,4,14), 151 => (2,4,14), 152 => (2,4,14), 153 => (2,4,14), 154 => (2,4,14), 155 => (2,4,14), 156 => (2,4,14), 157 => (2,4,14), 158 => (2,4,14), 159 => (2,4,14)), 
			77 => (0 => (2,4,14), 1 => (2,4,14), 2 => (2,4,14), 3 => (2,4,14), 4 => (2,4,14), 5 => (2,4,14), 6 => (2,4,14), 7 => (2,4,14), 8 => (2,4,14), 9 => (2,4,14), 10 => (2,4,14), 11 => (2,4,14), 12 => (2,4,14), 13 => (2,4,14), 14 => (2,4,14), 15 => (2,4,14), 16 => (2,4,14), 17 => (2,4,14), 18 => (2,4,14), 19 => (2,4,14), 20 => (2,4,14), 21 => (2,4,14), 22 => (2,4,14), 23 => (2,4,14), 24 => (2,4,14), 25 => (2,4,14), 26 => (2,4,14), 27 => (2,4,14), 28 => (0,4,15), 29 => (11,3,4), 30 => (14,15,15), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,12,7), 38 => (14,10,0), 39 => (12,8,0), 40 => (10,6,0), 41 => (5,0,0), 42 => (0,0,0), 43 => (1,0,0), 44 => (1,0,0), 45 => (3,1,0), 46 => (10,0,0), 47 => (1,4,15), 48 => (2,4,14), 49 => (2,4,14), 50 => (2,4,14), 51 => (2,4,14), 52 => (2,4,14), 53 => (2,4,14), 54 => (2,4,14), 55 => (2,4,14), 56 => (2,4,14), 57 => (2,4,14), 58 => (2,4,14), 59 => (2,4,14), 60 => (2,4,15), 61 => (0,0,3), 62 => (4,4,10), 63 => (7,7,15), 64 => (0,1,13), 65 => (4,4,15), 66 => (13,13,7), 67 => (15,15,0), 68 => (14,14,0), 69 => (14,14,0), 70 => (14,14,0), 71 => (15,15,3), 72 => (1,1,6), 73 => (2,2,10), 74 => (7,7,15), 75 => (10,10,14), 76 => (9,9,14), 77 => (12,12,14), 78 => (14,14,14), 79 => (15,15,14), 80 => (15,15,14), 81 => (15,15,14), 82 => (15,15,14), 83 => (9,9,14), 84 => (7,7,14), 85 => (5,5,15), 86 => (2,2,10), 87 => (2,2,6), 88 => (15,15,3), 89 => (14,14,0), 90 => (14,14,0), 91 => (14,14,0), 92 => (15,15,0), 93 => (13,13,7), 94 => (4,4,15), 95 => (0,1,13), 96 => (7,7,15), 97 => (4,4,10), 98 => (0,0,3), 99 => (2,4,15), 100 => (2,4,14), 101 => (2,4,14), 102 => (2,4,14), 103 => (2,4,14), 104 => (2,4,14), 105 => (2,4,14), 106 => (2,4,14), 107 => (2,4,14), 108 => (2,4,14), 109 => (2,4,14), 110 => (2,4,14), 111 => (2,4,14), 112 => (1,4,15), 113 => (10,0,0), 114 => (3,1,0), 115 => (1,0,0), 116 => (1,0,0), 117 => (0,0,0), 118 => (5,0,0), 119 => (10,6,0), 120 => (12,8,0), 121 => (14,10,0), 122 => (14,12,7), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,15,15), 130 => (11,3,4), 131 => (0,4,15), 132 => (2,4,14), 133 => (2,4,14), 134 => (2,4,14), 135 => (2,4,14), 136 => (2,4,14), 137 => (2,4,14), 138 => (2,4,14), 139 => (2,4,14), 140 => (2,4,14), 141 => (2,4,14), 142 => (2,4,14), 143 => (2,4,14), 144 => (2,4,14), 145 => (2,4,14), 146 => (2,4,14), 147 => (2,4,14), 148 => (2,4,14), 149 => (2,4,14), 150 => (2,4,14), 151 => (2,4,14), 152 => (2,4,14), 153 => (2,4,14), 154 => (2,4,14), 155 => (2,4,14), 156 => (2,4,14), 157 => (2,4,14), 158 => (2,4,14), 159 => (2,4,14)), 
			78 => (0 => (2,4,14), 1 => (2,4,14), 2 => (2,4,14), 3 => (2,4,14), 4 => (2,4,14), 5 => (2,4,14), 6 => (2,4,14), 7 => (2,4,14), 8 => (2,4,14), 9 => (2,4,14), 10 => (2,4,14), 11 => (2,4,14), 12 => (2,4,14), 13 => (2,4,14), 14 => (2,4,14), 15 => (2,4,14), 16 => (2,4,14), 17 => (2,4,14), 18 => (2,4,14), 19 => (2,4,14), 20 => (2,4,14), 21 => (2,4,14), 22 => (2,4,14), 23 => (2,4,14), 24 => (2,4,14), 25 => (2,4,14), 26 => (2,4,14), 27 => (2,4,14), 28 => (2,4,14), 29 => (0,3,15), 30 => (14,5,3), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,12,7), 38 => (14,10,0), 39 => (12,8,0), 40 => (10,6,0), 41 => (9,3,0), 42 => (7,0,0), 43 => (4,0,0), 44 => (1,0,0), 45 => (3,1,0), 46 => (10,0,0), 47 => (1,4,15), 48 => (2,4,14), 49 => (2,4,14), 50 => (2,4,14), 51 => (2,4,14), 52 => (2,4,14), 53 => (2,4,14), 54 => (2,4,14), 55 => (2,4,14), 56 => (2,4,14), 57 => (2,4,14), 58 => (2,4,14), 59 => (2,4,14), 60 => (2,4,14), 61 => (2,4,15), 62 => (1,2,10), 63 => (0,0,4), 64 => (6,6,14), 65 => (7,7,14), 66 => (3,3,14), 67 => (5,5,15), 68 => (13,13,6), 69 => (13,13,2), 70 => (15,15,0), 71 => (7,7,7), 72 => (0,0,13), 73 => (0,0,12), 74 => (1,1,13), 75 => (5,5,14), 76 => (6,6,14), 77 => (6,6,14), 78 => (8,8,14), 79 => (12,12,14), 80 => (12,12,14), 81 => (12,12,14), 82 => (13,13,14), 83 => (10,10,14), 84 => (4,4,14), 85 => (2,2,13), 86 => (0,0,11), 87 => (0,0,14), 88 => (3,3,7), 89 => (15,15,0), 90 => (13,13,2), 91 => (13,13,6), 92 => (5,5,15), 93 => (3,3,14), 94 => (7,7,14), 95 => (6,6,14), 96 => (0,0,4), 97 => (1,2,10), 98 => (2,4,15), 99 => (2,4,14), 100 => (2,4,14), 101 => (2,4,14), 102 => (2,4,14), 103 => (2,4,14), 104 => (2,4,14), 105 => (2,4,14), 106 => (2,4,14), 107 => (2,4,14), 108 => (2,4,14), 109 => (2,4,14), 110 => (2,4,14), 111 => (2,4,14), 112 => (1,4,15), 113 => (10,0,0), 114 => (3,1,0), 115 => (1,0,0), 116 => (4,0,0), 117 => (7,0,0), 118 => (9,3,0), 119 => (10,6,0), 120 => (12,8,0), 121 => (14,10,0), 122 => (14,12,7), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,5,3), 130 => (0,3,15), 131 => (2,4,14), 132 => (2,4,14), 133 => (2,4,14), 134 => (2,4,14), 135 => (2,4,14), 136 => (2,4,14), 137 => (2,4,14), 138 => (2,4,14), 139 => (2,4,14), 140 => (2,4,14), 141 => (2,4,14), 142 => (2,4,14), 143 => (2,4,14), 144 => (2,4,14), 145 => (2,4,14), 146 => (2,4,14), 147 => (2,4,14), 148 => (2,4,14), 149 => (2,4,14), 150 => (2,4,14), 151 => (2,4,14), 152 => (2,4,14), 153 => (2,4,14), 154 => (2,4,14), 155 => (2,4,14), 156 => (2,4,14), 157 => (2,4,14), 158 => (2,4,14), 159 => (2,4,14)), 
			79 => (0 => (1,3,14), 1 => (1,3,14), 2 => (1,3,14), 3 => (1,3,14), 4 => (1,3,14), 5 => (1,3,14), 6 => (1,3,14), 7 => (1,3,14), 8 => (1,3,14), 9 => (1,3,14), 10 => (1,3,14), 11 => (1,3,14), 12 => (1,3,14), 13 => (1,3,14), 14 => (1,3,14), 15 => (1,3,14), 16 => (1,3,14), 17 => (1,3,14), 18 => (1,3,14), 19 => (1,3,14), 20 => (1,3,14), 21 => (1,3,14), 22 => (1,3,14), 23 => (1,3,14), 24 => (1,3,14), 25 => (1,3,14), 26 => (1,3,14), 27 => (1,3,14), 28 => (1,4,14), 29 => (3,1,10), 30 => (14,11,10), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,14,14), 37 => (14,12,7), 38 => (14,10,0), 39 => (12,9,0), 40 => (9,4,0), 41 => (4,1,0), 42 => (0,0,0), 43 => (5,0,0), 44 => (3,0,0), 45 => (3,0,0), 46 => (9,0,0), 47 => (1,4,15), 48 => (1,3,14), 49 => (1,3,14), 50 => (1,3,14), 51 => (1,3,14), 52 => (1,3,14), 53 => (1,3,14), 54 => (1,3,14), 55 => (1,3,14), 56 => (1,3,14), 57 => (1,3,14), 58 => (1,3,14), 59 => (1,3,14), 60 => (1,3,14), 61 => (1,3,14), 62 => (1,4,14), 63 => (2,4,15), 64 => (0,2,9), 65 => (1,2,8), 66 => (6,6,14), 67 => (7,7,14), 68 => (3,3,15), 69 => (4,4,15), 70 => (11,11,15), 71 => (0,0,4), 72 => (0,0,12), 73 => (0,0,12), 74 => (0,0,11), 75 => (0,0,11), 76 => (0,0,12), 77 => (4,4,14), 78 => (8,8,14), 79 => (7,7,14), 80 => (7,7,14), 81 => (7,7,14), 82 => (8,8,14), 83 => (13,13,14), 84 => (7,7,14), 85 => (1,1,12), 86 => (0,0,11), 87 => (0,0,12), 88 => (0,0,4), 89 => (9,9,15), 90 => (4,4,15), 91 => (3,3,15), 92 => (7,7,14), 93 => (6,6,14), 94 => (1,2,8), 95 => (0,2,9), 96 => (2,4,15), 97 => (1,4,14), 98 => (1,3,14), 99 => (1,3,14), 100 => (1,3,14), 101 => (1,3,14), 102 => (1,3,14), 103 => (1,3,14), 104 => (1,3,14), 105 => (1,3,14), 106 => (1,3,14), 107 => (1,3,14), 108 => (1,3,14), 109 => (1,3,14), 110 => (1,3,14), 111 => (1,3,14), 112 => (1,4,15), 113 => (9,0,0), 114 => (3,0,0), 115 => (3,0,0), 116 => (5,0,0), 117 => (0,0,0), 118 => (4,1,0), 119 => (9,4,0), 120 => (12,9,0), 121 => (14,10,0), 122 => (14,12,7), 123 => (14,14,14), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,11,10), 130 => (3,1,10), 131 => (1,4,14), 132 => (1,3,14), 133 => (1,3,14), 134 => (1,3,14), 135 => (1,3,14), 136 => (1,3,14), 137 => (1,3,14), 138 => (1,3,14), 139 => (1,3,14), 140 => (1,3,14), 141 => (1,3,14), 142 => (1,3,14), 143 => (1,3,14), 144 => (1,3,14), 145 => (1,3,14), 146 => (1,3,14), 147 => (1,3,14), 148 => (1,3,14), 149 => (1,3,14), 150 => (1,3,14), 151 => (1,3,14), 152 => (1,3,14), 153 => (1,3,14), 154 => (1,3,14), 155 => (1,3,14), 156 => (1,3,14), 157 => (1,3,14), 158 => (1,3,14), 159 => (1,3,14)), 
			80 => (0 => (3,5,14), 1 => (3,5,14), 2 => (3,5,14), 3 => (3,5,14), 4 => (3,5,14), 5 => (3,5,14), 6 => (3,5,14), 7 => (3,5,14), 8 => (3,5,14), 9 => (3,5,14), 10 => (3,5,14), 11 => (3,5,14), 12 => (3,5,14), 13 => (3,5,14), 14 => (3,5,14), 15 => (3,5,14), 16 => (3,5,14), 17 => (3,5,14), 18 => (3,5,14), 19 => (3,5,14), 20 => (3,5,14), 21 => (3,5,14), 22 => (3,5,14), 23 => (3,5,14), 24 => (3,5,14), 25 => (3,5,14), 26 => (3,5,14), 27 => (3,5,14), 28 => (1,5,15), 29 => (11,3,4), 30 => (14,15,15), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,14,14), 34 => (14,14,14), 35 => (14,14,14), 36 => (14,15,15), 37 => (15,14,7), 38 => (9,4,0), 39 => (6,0,0), 40 => (5,0,0), 41 => (3,0,0), 42 => (1,0,0), 43 => (1,0,0), 44 => (2,0,0), 45 => (0,0,0), 46 => (6,0,0), 47 => (2,5,15), 48 => (3,5,14), 49 => (3,5,14), 50 => (3,5,14), 51 => (3,5,14), 52 => (3,5,14), 53 => (3,5,14), 54 => (3,5,14), 55 => (3,5,14), 56 => (3,5,14), 57 => (3,5,14), 58 => (3,5,14), 59 => (3,5,14), 60 => (3,5,14), 61 => (3,5,14), 62 => (3,5,14), 63 => (3,5,14), 64 => (3,5,14), 65 => (3,5,15), 66 => (0,1,4), 67 => (1,2,9), 68 => (3,3,8), 69 => (7,7,15), 70 => (12,12,15), 71 => (0,0,4), 72 => (0,0,12), 73 => (0,0,12), 74 => (0,0,12), 75 => (0,0,11), 76 => (0,0,12), 77 => (5,5,15), 78 => (10,10,14), 79 => (6,6,14), 80 => (4,4,14), 81 => (4,4,14), 82 => (4,4,14), 83 => (6,6,14), 84 => (10,10,14), 85 => (1,1,12), 86 => (0,0,11), 87 => (0,0,12), 88 => (0,0,4), 89 => (10,10,15), 90 => (8,7,15), 91 => (3,3,8), 92 => (2,3,9), 93 => (0,1,4), 94 => (3,5,15), 95 => (3,5,14), 96 => (3,5,14), 97 => (3,5,14), 98 => (3,5,14), 99 => (3,5,14), 100 => (3,5,14), 101 => (3,5,14), 102 => (3,5,14), 103 => (3,5,14), 104 => (3,5,14), 105 => (3,5,14), 106 => (3,5,14), 107 => (3,5,14), 108 => (3,5,14), 109 => (3,5,14), 110 => (3,5,14), 111 => (3,5,14), 112 => (2,5,15), 113 => (6,0,0), 114 => (0,0,0), 115 => (2,0,0), 116 => (1,0,0), 117 => (1,0,0), 118 => (3,0,0), 119 => (5,0,0), 120 => (6,0,0), 121 => (9,4,0), 122 => (15,14,7), 123 => (14,15,15), 124 => (14,14,14), 125 => (14,14,14), 126 => (14,14,14), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,15,15), 130 => (10,2,4), 131 => (1,5,15), 132 => (3,5,14), 133 => (3,5,14), 134 => (3,5,14), 135 => (3,5,14), 136 => (3,5,14), 137 => (3,5,14), 138 => (3,5,14), 139 => (3,5,14), 140 => (3,5,14), 141 => (3,5,14), 142 => (3,5,14), 143 => (3,5,14), 144 => (3,5,14), 145 => (3,5,14), 146 => (3,5,14), 147 => (3,5,14), 148 => (3,5,14), 149 => (3,5,14), 150 => (3,5,14), 151 => (3,5,14), 152 => (3,5,14), 153 => (3,5,14), 154 => (3,5,14), 155 => (3,5,14), 156 => (3,5,14), 157 => (3,5,14), 158 => (3,5,14), 159 => (3,5,14)), 
			81 => (0 => (3,5,14), 1 => (3,5,14), 2 => (3,5,14), 3 => (3,5,14), 4 => (3,5,14), 5 => (3,5,14), 6 => (3,5,14), 7 => (3,5,14), 8 => (3,5,14), 9 => (3,5,14), 10 => (3,5,14), 11 => (3,5,14), 12 => (3,5,14), 13 => (3,5,14), 14 => (3,5,14), 15 => (3,5,14), 16 => (3,5,14), 17 => (3,5,14), 18 => (3,5,14), 19 => (3,5,14), 20 => (3,5,14), 21 => (3,5,14), 22 => (3,5,14), 23 => (3,5,14), 24 => (3,5,14), 25 => (3,5,14), 26 => (3,5,14), 27 => (2,5,14), 28 => (3,2,10), 29 => (14,11,10), 30 => (14,14,14), 31 => (14,14,14), 32 => (14,14,14), 33 => (14,15,15), 34 => (14,15,15), 35 => (12,6,6), 36 => (12,2,2), 37 => (8,0,0), 38 => (5,0,0), 39 => (5,0,0), 40 => (6,0,0), 41 => (4,0,0), 42 => (1,0,0), 43 => (2,0,0), 44 => (1,0,0), 45 => (0,0,0), 46 => (9,2,7), 47 => (2,5,14), 48 => (3,5,14), 49 => (3,5,14), 50 => (3,5,14), 51 => (3,5,14), 52 => (3,5,14), 53 => (3,5,14), 54 => (3,5,14), 55 => (3,5,14), 56 => (3,5,14), 57 => (3,5,14), 58 => (3,5,14), 59 => (3,5,14), 60 => (3,5,14), 61 => (3,5,14), 62 => (3,5,14), 63 => (3,5,14), 64 => (3,5,14), 65 => (3,5,14), 66 => (3,5,14), 67 => (3,5,14), 68 => (3,5,15), 69 => (0,0,4), 70 => (8,8,10), 71 => (0,0,4), 72 => (0,0,12), 73 => (0,0,11), 74 => (0,0,11), 75 => (2,2,13), 76 => (6,6,6), 77 => (7,7,7), 78 => (6,6,7), 79 => (5,5,7), 80 => (5,5,7), 81 => (5,5,7), 82 => (5,5,7), 83 => (6,6,6), 84 => (7,7,14), 85 => (6,6,13), 86 => (0,0,11), 87 => (0,0,12), 88 => (0,0,4), 89 => (5,5,10), 90 => (0,1,4), 91 => (3,5,15), 92 => (3,5,14), 93 => (3,5,14), 94 => (3,5,14), 95 => (3,5,14), 96 => (3,5,14), 97 => (3,5,14), 98 => (3,5,14), 99 => (3,5,14), 100 => (3,5,14), 101 => (3,5,14), 102 => (3,5,14), 103 => (3,5,14), 104 => (3,5,14), 105 => (3,5,14), 106 => (3,5,14), 107 => (3,5,14), 108 => (3,5,14), 109 => (3,5,14), 110 => (3,5,14), 111 => (3,5,14), 112 => (2,5,14), 113 => (9,2,7), 114 => (0,0,0), 115 => (1,0,0), 116 => (2,0,0), 117 => (1,0,0), 118 => (4,0,0), 119 => (6,0,0), 120 => (5,0,0), 121 => (5,0,0), 122 => (8,0,0), 123 => (12,2,2), 124 => (12,6,6), 125 => (14,15,15), 126 => (14,15,15), 127 => (14,14,14), 128 => (14,14,14), 129 => (14,14,14), 130 => (14,11,10), 131 => (4,2,10), 132 => (2,5,14), 133 => (3,5,14), 134 => (3,5,14), 135 => (3,5,14), 136 => (3,5,14), 137 => (3,5,14), 138 => (3,5,14), 139 => (3,5,14), 140 => (3,5,14), 141 => (3,5,14), 142 => (3,5,14), 143 => (3,5,14), 144 => (3,5,14), 145 => (3,5,14), 146 => (3,5,14), 147 => (3,5,14), 148 => (3,5,14), 149 => (3,5,14), 150 => (3,5,14), 151 => (3,5,14), 152 => (3,5,14), 153 => (3,5,14), 154 => (3,5,14), 155 => (3,5,14), 156 => (3,5,14), 157 => (3,5,14), 158 => (3,5,14), 159 => (3,5,14)), 
			82 => (0 => (2,4,14), 1 => (2,4,14), 2 => (2,4,14), 3 => (2,4,14), 4 => (2,4,14), 5 => (2,4,14), 6 => (2,4,14), 7 => (2,4,14), 8 => (2,4,14), 9 => (2,4,14), 10 => (2,4,14), 11 => (2,4,14), 12 => (2,4,14), 13 => (2,4,14), 14 => (2,4,14), 15 => (2,4,14), 16 => (2,4,14), 17 => (2,4,14), 18 => (2,4,14), 19 => (2,4,14), 20 => (2,4,14), 21 => (2,4,14), 22 => (2,4,14), 23 => (2,4,14), 24 => (2,4,14), 25 => (2,4,14), 26 => (2,4,14), 27 => (1,5,15), 28 => (11,4,5), 29 => (14,15,15), 30 => (14,15,15), 31 => (13,11,11), 32 => (13,7,7), 33 => (12,2,2), 34 => (11,0,0), 35 => (11,0,0), 36 => (12,0,0), 37 => (9,0,0), 38 => (5,0,0), 39 => (6,0,0), 40 => (6,0,0), 41 => (4,0,0), 42 => (1,0,0), 43 => (1,0,0), 44 => (4,0,0), 45 => (9,0,1), 46 => (1,5,15), 47 => (2,4,14), 48 => (2,4,14), 49 => (2,4,14), 50 => (2,4,14), 51 => (2,4,14), 52 => (2,4,14), 53 => (2,4,14), 54 => (2,4,14), 55 => (2,4,14), 56 => (2,4,14), 57 => (2,4,14), 58 => (2,4,14), 59 => (2,4,14), 60 => (2,4,14), 61 => (2,4,14), 62 => (2,4,14), 63 => (2,4,14), 64 => (2,4,14), 65 => (2,4,14), 66 => (2,4,14), 67 => (2,4,14), 68 => (2,4,14), 69 => (2,5,15), 70 => (8,8,5), 71 => (6,6,11), 72 => (6,6,15), 73 => (6,6,14), 74 => (5,5,14), 75 => (9,9,15), 76 => (0,0,0), 77 => (0,0,0), 78 => (0,0,0), 79 => (0,0,0), 80 => (0,0,0), 81 => (0,0,0), 82 => (0,0,0), 83 => (0,0,0), 84 => (5,5,14), 85 => (0,0,12), 86 => (4,4,13), 87 => (0,0,12), 88 => (0,0,5), 89 => (5,5,5), 90 => (2,5,15), 91 => (2,4,14), 92 => (2,4,14), 93 => (2,4,14), 94 => (2,4,14), 95 => (2,4,14), 96 => (2,4,14), 97 => (2,4,14), 98 => (2,4,14), 99 => (2,4,14), 100 => (2,4,14), 101 => (2,4,14), 102 => (2,4,14), 103 => (2,4,14), 104 => (2,4,14), 105 => (2,4,14), 106 => (2,4,14), 107 => (2,4,14), 108 => (2,4,14), 109 => (2,4,14), 110 => (2,4,14), 111 => (2,4,14), 112 => (2,4,14), 113 => (1,5,15), 114 => (9,0,1), 115 => (4,0,0), 116 => (1,0,0), 117 => (1,0,0), 118 => (4,0,0), 119 => (6,0,0), 120 => (6,0,0), 121 => (5,0,0), 122 => (9,0,0), 123 => (12,0,0), 124 => (11,0,0), 125 => (11,0,0), 126 => (12,2,2), 127 => (13,7,7), 128 => (13,11,11), 129 => (14,15,15), 130 => (14,15,15), 131 => (10,3,5), 132 => (1,5,15), 133 => (2,4,14), 134 => (2,4,14), 135 => (2,4,14), 136 => (2,4,14), 137 => (2,4,14), 138 => (2,4,14), 139 => (2,4,14), 140 => (2,4,14), 141 => (2,4,14), 142 => (2,4,14), 143 => (2,4,14), 144 => (2,4,14), 145 => (2,4,14), 146 => (2,4,14), 147 => (2,4,14), 148 => (2,4,14), 149 => (2,4,14), 150 => (2,4,14), 151 => (2,4,14), 152 => (2,4,14), 153 => (2,4,14), 154 => (2,4,14), 155 => (2,4,14), 156 => (2,4,14), 157 => (2,4,14), 158 => (2,4,14), 159 => (2,4,14)), 
			83 => (0 => (3,5,14), 1 => (3,5,14), 2 => (3,5,14), 3 => (3,5,14), 4 => (3,5,14), 5 => (3,5,14), 6 => (3,5,14), 7 => (3,5,14), 8 => (3,5,14), 9 => (3,5,14), 10 => (3,5,14), 11 => (3,5,14), 12 => (3,5,14), 13 => (3,5,14), 14 => (3,5,14), 15 => (3,5,14), 16 => (3,5,14), 17 => (3,5,14), 18 => (3,5,14), 19 => (3,5,14), 20 => (3,5,14), 21 => (3,5,14), 22 => (3,5,14), 23 => (3,5,14), 24 => (3,5,14), 25 => (3,5,14), 26 => (3,5,14), 27 => (4,4,11), 28 => (13,3,2), 29 => (12,3,3), 30 => (11,0,0), 31 => (11,0,0), 32 => (11,0,0), 33 => (11,0,0), 34 => (12,0,0), 35 => (12,0,0), 36 => (12,0,0), 37 => (9,0,0), 38 => (5,0,0), 39 => (6,0,0), 40 => (6,0,0), 41 => (3,0,0), 42 => (4,0,0), 43 => (9,1,2), 44 => (5,4,11), 45 => (2,6,15), 46 => (3,5,14), 47 => (3,5,14), 48 => (3,5,14), 49 => (3,5,14), 50 => (3,5,14), 51 => (3,5,14), 52 => (3,5,14), 53 => (3,5,14), 54 => (3,5,14), 55 => (3,5,14), 56 => (3,5,14), 57 => (3,5,14), 58 => (3,5,14), 59 => (3,5,14), 60 => (3,5,14), 61 => (3,5,14), 62 => (3,5,14), 63 => (3,5,14), 64 => (3,5,14), 65 => (3,5,14), 66 => (3,5,14), 67 => (3,5,14), 68 => (3,5,14), 69 => (3,5,14), 70 => (1,2,6), 71 => (0,0,0), 72 => (0,0,0), 73 => (0,0,0), 74 => (2,2,1), 75 => (5,5,6), 76 => (9,9,7), 77 => (5,5,7), 78 => (8,9,15), 79 => (8,9,15), 80 => (7,10,13), 81 => (5,11,9), 82 => (10,14,7), 83 => (5,5,7), 84 => (6,6,14), 85 => (0,0,11), 86 => (1,1,12), 87 => (1,1,13), 88 => (0,0,4), 89 => (7,8,15), 90 => (3,5,14), 91 => (3,5,14), 92 => (3,5,14), 93 => (3,5,14), 94 => (3,5,14), 95 => (3,5,14), 96 => (3,5,14), 97 => (3,5,14), 98 => (3,5,14), 99 => (3,5,14), 100 => (3,5,14), 101 => (3,5,14), 102 => (3,5,14), 103 => (3,5,14), 104 => (3,5,14), 105 => (3,5,14), 106 => (3,5,14), 107 => (3,5,14), 108 => (3,5,14), 109 => (3,5,14), 110 => (3,5,14), 111 => (3,5,14), 112 => (3,5,14), 113 => (3,5,14), 114 => (2,6,15), 115 => (6,5,11), 116 => (9,0,2), 117 => (4,0,0), 118 => (3,0,0), 119 => (6,0,0), 120 => (6,0,0), 121 => (5,0,0), 122 => (9,0,0), 123 => (12,0,0), 124 => (12,0,0), 125 => (12,0,0), 126 => (11,0,0), 127 => (11,0,0), 128 => (11,0,0), 129 => (11,0,0), 130 => (12,3,3), 131 => (13,3,2), 132 => (4,4,11), 133 => (3,5,14), 134 => (3,5,14), 135 => (3,5,14), 136 => (3,5,14), 137 => (3,5,14), 138 => (3,5,14), 139 => (3,5,14), 140 => (3,5,14), 141 => (3,5,14), 142 => (3,5,14), 143 => (3,5,14), 144 => (3,5,14), 145 => (3,5,14), 146 => (3,5,14), 147 => (3,5,14), 148 => (3,5,14), 149 => (3,5,14), 150 => (3,5,14), 151 => (3,5,14), 152 => (3,5,14), 153 => (3,5,14), 154 => (3,5,14), 155 => (3,5,14), 156 => (3,5,14), 157 => (3,5,14), 158 => (3,5,14), 159 => (3,5,14)), 
			84 => (0 => (3,5,14), 1 => (3,5,14), 2 => (3,5,14), 3 => (3,5,14), 4 => (3,5,14), 5 => (3,5,14), 6 => (3,5,14), 7 => (3,5,14), 8 => (3,5,14), 9 => (3,5,14), 10 => (3,5,14), 11 => (3,5,14), 12 => (3,5,14), 13 => (3,5,14), 14 => (3,5,14), 15 => (3,5,14), 16 => (3,5,14), 17 => (3,5,14), 18 => (3,5,14), 19 => (3,5,14), 20 => (3,5,14), 21 => (3,5,14), 22 => (3,5,14), 23 => (3,5,14), 24 => (3,5,14), 25 => (3,5,14), 26 => (2,6,15), 27 => (10,1,2), 28 => (12,0,0), 29 => (11,0,0), 30 => (12,0,0), 31 => (12,0,0), 32 => (12,0,0), 33 => (12,0,0), 34 => (12,0,0), 35 => (12,0,0), 36 => (12,0,0), 37 => (8,0,0), 38 => (5,0,0), 39 => (5,0,0), 40 => (7,0,0), 41 => (9,0,2), 42 => (6,4,11), 43 => (3,6,15), 44 => (3,6,14), 45 => (3,5,14), 46 => (3,5,14), 47 => (3,5,14), 48 => (3,5,14), 49 => (3,5,14), 50 => (3,5,14), 51 => (3,5,14), 52 => (3,5,14), 53 => (3,5,14), 54 => (3,5,14), 55 => (3,5,14), 56 => (3,5,14), 57 => (3,5,14), 58 => (3,5,14), 59 => (3,5,14), 60 => (3,5,14), 61 => (3,5,14), 62 => (3,5,14), 63 => (3,5,14), 64 => (3,5,14), 65 => (3,5,14), 66 => (3,5,14), 67 => (3,5,14), 68 => (3,5,14), 69 => (3,5,14), 70 => (4,6,15), 71 => (1,2,6), 72 => (3,3,2), 73 => (9,9,8), 74 => (2,2,6), 75 => (0,0,4), 76 => (1,1,5), 77 => (0,0,5), 78 => (0,0,4), 79 => (0,0,4), 80 => (0,0,4), 81 => (0,0,5), 82 => (0,0,5), 83 => (0,0,4), 84 => (0,0,8), 85 => (0,0,12), 86 => (0,0,11), 87 => (0,0,12), 88 => (0,0,4), 89 => (8,9,15), 90 => (3,5,14), 91 => (3,5,14), 92 => (3,5,14), 93 => (3,5,14), 94 => (3,5,14), 95 => (3,5,14), 96 => (3,5,14), 97 => (3,5,14), 98 => (3,5,14), 99 => (3,5,14), 100 => (3,5,14), 101 => (3,5,14), 102 => (3,5,14), 103 => (3,5,14), 104 => (3,5,14), 105 => (3,5,14), 106 => (3,5,14), 107 => (3,5,14), 108 => (3,5,14), 109 => (3,5,14), 110 => (3,5,14), 111 => (3,5,14), 112 => (3,5,14), 113 => (3,5,14), 114 => (3,5,14), 115 => (3,5,14), 116 => (3,6,15), 117 => (6,4,11), 118 => (9,0,2), 119 => (7,0,0), 120 => (5,0,0), 121 => (5,0,0), 122 => (8,0,0), 123 => (12,0,0), 124 => (12,0,0), 125 => (12,0,0), 126 => (12,0,0), 127 => (12,0,0), 128 => (12,0,0), 129 => (12,0,0), 130 => (11,0,0), 131 => (12,0,0), 132 => (10,1,2), 133 => (3,6,15), 134 => (3,5,14), 135 => (3,5,14), 136 => (3,5,14), 137 => (3,5,14), 138 => (3,5,14), 139 => (3,5,14), 140 => (3,5,14), 141 => (3,5,14), 142 => (3,5,14), 143 => (3,5,14), 144 => (3,5,14), 145 => (3,5,14), 146 => (3,5,14), 147 => (3,5,14), 148 => (3,5,14), 149 => (3,5,14), 150 => (3,5,14), 151 => (3,5,14), 152 => (3,5,14), 153 => (3,5,14), 154 => (3,5,14), 155 => (3,5,14), 156 => (3,5,14), 157 => (3,5,14), 158 => (3,5,14), 159 => (3,5,14)), 
			85 => (0 => (5,8,14), 1 => (5,8,14), 2 => (5,8,14), 3 => (5,8,14), 4 => (5,8,14), 5 => (5,8,14), 6 => (5,8,14), 7 => (5,8,14), 8 => (5,8,14), 9 => (5,8,14), 10 => (5,8,14), 11 => (5,8,14), 12 => (5,8,14), 13 => (5,8,14), 14 => (5,8,14), 15 => (5,8,14), 16 => (5,8,14), 17 => (5,8,14), 18 => (5,8,14), 19 => (5,8,14), 20 => (5,8,14), 21 => (5,8,14), 22 => (5,8,14), 23 => (5,8,14), 24 => (5,8,14), 25 => (4,8,14), 26 => (6,7,11), 27 => (12,0,0), 28 => (12,0,0), 29 => (12,0,0), 30 => (12,0,0), 31 => (12,0,0), 32 => (12,0,0), 33 => (12,0,0), 34 => (12,0,0), 35 => (12,0,0), 36 => (12,0,0), 37 => (11,0,0), 38 => (9,0,0), 39 => (9,4,7), 40 => (7,7,11), 41 => (4,9,15), 42 => (4,8,14), 43 => (5,8,14), 44 => (5,8,14), 45 => (5,8,14), 46 => (5,8,14), 47 => (5,8,14), 48 => (5,8,14), 49 => (5,8,14), 50 => (5,8,14), 51 => (5,8,14), 52 => (5,8,14), 53 => (5,8,14), 54 => (5,8,14), 55 => (5,8,14), 56 => (5,8,14), 57 => (5,8,14), 58 => (5,8,14), 59 => (5,8,14), 60 => (5,8,14), 61 => (5,8,14), 62 => (5,8,14), 63 => (5,8,14), 64 => (5,8,14), 65 => (5,8,14), 66 => (5,8,14), 67 => (5,8,14), 68 => (5,8,14), 69 => (5,8,14), 70 => (4,8,14), 71 => (8,12,15), 72 => (3,3,5), 73 => (0,0,8), 74 => (0,0,13), 75 => (1,1,13), 76 => (2,2,13), 77 => (0,0,12), 78 => (0,0,12), 79 => (0,0,12), 80 => (0,0,12), 81 => (0,0,12), 82 => (0,0,12), 83 => (0,0,12), 84 => (0,0,12), 85 => (0,0,12), 86 => (0,0,12), 87 => (0,0,12), 88 => (0,0,3), 89 => (8,10,15), 90 => (4,7,14), 91 => (5,8,14), 92 => (5,8,14), 93 => (5,8,14), 94 => (5,8,14), 95 => (5,8,14), 96 => (5,8,14), 97 => (5,8,14), 98 => (5,8,14), 99 => (5,8,14), 100 => (5,8,14), 101 => (5,8,14), 102 => (5,8,14), 103 => (5,8,14), 104 => (5,8,14), 105 => (5,8,14), 106 => (5,8,14), 107 => (5,8,14), 108 => (5,8,14), 109 => (5,8,14), 110 => (5,8,14), 111 => (5,8,14), 112 => (5,8,14), 113 => (5,8,14), 114 => (5,8,14), 115 => (5,8,14), 116 => (5,8,14), 117 => (4,8,14), 118 => (4,9,15), 119 => (6,5,11), 120 => (9,4,7), 121 => (9,0,0), 122 => (11,0,0), 123 => (12,0,0), 124 => (12,0,0), 125 => (12,0,0), 126 => (12,0,0), 127 => (12,0,0), 128 => (12,0,0), 129 => (12,0,0), 130 => (12,0,0), 131 => (12,0,0), 132 => (12,0,0), 133 => (5,6,11), 134 => (4,8,14), 135 => (5,8,14), 136 => (5,8,14), 137 => (5,8,14), 138 => (5,8,14), 139 => (5,8,14), 140 => (5,8,14), 141 => (5,8,14), 142 => (5,8,14), 143 => (5,8,14), 144 => (5,8,14), 145 => (5,8,14), 146 => (5,8,14), 147 => (5,8,14), 148 => (5,8,14), 149 => (5,8,14), 150 => (5,8,14), 151 => (5,8,14), 152 => (5,8,14), 153 => (5,8,14), 154 => (5,8,14), 155 => (5,8,14), 156 => (5,8,14), 157 => (5,8,14), 158 => (5,8,14), 159 => (5,8,14)), 
			86 => (0 => (4,7,14), 1 => (4,7,14), 2 => (4,7,14), 3 => (4,7,14), 4 => (4,7,14), 5 => (4,7,14), 6 => (4,7,14), 7 => (4,7,14), 8 => (4,7,14), 9 => (4,7,14), 10 => (4,7,14), 11 => (4,7,14), 12 => (4,7,14), 13 => (4,7,14), 14 => (4,7,14), 15 => (4,7,14), 16 => (4,7,14), 17 => (4,7,14), 18 => (4,7,14), 19 => (4,7,14), 20 => (4,7,14), 21 => (4,7,14), 22 => (4,7,14), 23 => (4,7,14), 24 => (4,7,14), 25 => (4,8,15), 26 => (10,0,2), 27 => (12,0,0), 28 => (12,0,0), 29 => (12,0,0), 30 => (12,0,0), 31 => (12,0,0), 32 => (12,0,0), 33 => (12,0,0), 34 => (12,0,0), 35 => (13,0,0), 36 => (8,3,7), 37 => (6,7,11), 38 => (4,8,15), 39 => (4,8,14), 40 => (4,7,14), 41 => (4,7,14), 42 => (4,7,14), 43 => (4,7,14), 44 => (4,7,14), 45 => (4,7,14), 46 => (4,7,14), 47 => (4,7,14), 48 => (4,7,14), 49 => (4,7,14), 50 => (4,7,14), 51 => (4,7,14), 52 => (4,7,14), 53 => (4,7,14), 54 => (4,7,14), 55 => (4,7,14), 56 => (4,7,14), 57 => (4,7,14), 58 => (4,7,14), 59 => (4,7,14), 60 => (4,7,14), 61 => (4,7,14), 62 => (4,7,14), 63 => (4,7,14), 64 => (4,7,14), 65 => (4,7,14), 66 => (4,7,14), 67 => (4,7,14), 68 => (4,7,14), 69 => (4,7,14), 70 => (4,7,14), 71 => (9,9,9), 72 => (0,0,8), 73 => (0,0,12), 74 => (0,0,11), 75 => (4,4,13), 76 => (0,0,11), 77 => (0,0,12), 78 => (0,0,12), 79 => (0,0,12), 80 => (0,0,12), 81 => (0,0,12), 82 => (0,0,12), 83 => (0,0,12), 84 => (0,0,12), 85 => (0,0,12), 86 => (0,0,12), 87 => (0,0,12), 88 => (2,1,10), 89 => (8,10,1), 90 => (4,9,8), 91 => (1,7,7), 92 => (5,6,15), 93 => (5,8,15), 94 => (5,7,14), 95 => (4,7,14), 96 => (4,7,14), 97 => (4,7,14), 98 => (4,7,14), 99 => (4,7,14), 100 => (4,7,14), 101 => (4,7,14), 102 => (4,7,14), 103 => (4,7,14), 104 => (4,7,14), 105 => (4,7,14), 106 => (4,7,14), 107 => (4,7,14), 108 => (4,7,14), 109 => (4,7,14), 110 => (4,7,14), 111 => (4,7,14), 112 => (4,7,14), 113 => (4,7,14), 114 => (4,7,14), 115 => (4,7,14), 116 => (4,7,14), 117 => (4,7,14), 118 => (4,7,14), 119 => (4,8,14), 120 => (4,8,14), 121 => (4,9,15), 122 => (6,5,11), 123 => (8,4,7), 124 => (13,0,0), 125 => (12,0,0), 126 => (12,0,0), 127 => (12,0,0), 128 => (12,0,0), 129 => (12,0,0), 130 => (12,0,0), 131 => (12,0,0), 132 => (12,0,0), 133 => (11,2,2), 134 => (4,8,15), 135 => (4,7,14), 136 => (4,7,14), 137 => (4,7,14), 138 => (4,7,14), 139 => (4,7,14), 140 => (4,7,14), 141 => (4,7,14), 142 => (4,7,14), 143 => (4,7,14), 144 => (4,7,14), 145 => (4,7,14), 146 => (4,7,14), 147 => (4,7,14), 148 => (4,7,14), 149 => (4,7,14), 150 => (4,7,14), 151 => (4,7,14), 152 => (4,7,14), 153 => (4,7,14), 154 => (4,7,14), 155 => (4,7,14), 156 => (4,7,14), 157 => (4,7,14), 158 => (4,7,14), 159 => (4,7,14)), 
			87 => (0 => (6,10,14), 1 => (6,10,14), 2 => (6,10,14), 3 => (6,10,14), 4 => (6,10,14), 5 => (6,10,14), 6 => (6,10,14), 7 => (6,10,14), 8 => (6,10,14), 9 => (6,10,14), 10 => (6,10,14), 11 => (6,10,14), 12 => (6,10,14), 13 => (6,10,14), 14 => (6,10,14), 15 => (6,10,14), 16 => (6,10,14), 17 => (6,10,14), 18 => (6,10,14), 19 => (6,10,14), 20 => (6,10,14), 21 => (6,10,14), 22 => (6,10,14), 23 => (6,10,14), 24 => (5,10,14), 25 => (7,8,11), 26 => (12,0,0), 27 => (12,0,0), 28 => (12,0,0), 29 => (12,0,0), 30 => (12,0,0), 31 => (13,0,0), 32 => (8,5,7), 33 => (9,4,6), 34 => (4,11,15), 35 => (5,11,15), 36 => (5,10,14), 37 => (5,10,14), 38 => (6,10,14), 39 => (6,10,14), 40 => (6,10,14), 41 => (6,10,14), 42 => (6,10,14), 43 => (6,10,14), 44 => (6,10,15), 45 => (6,10,15), 46 => (6,10,15), 47 => (5,9,15), 48 => (6,10,15), 49 => (6,10,14), 50 => (6,10,14), 51 => (6,10,14), 52 => (6,10,14), 53 => (6,10,14), 54 => (6,10,14), 55 => (6,10,14), 56 => (6,10,14), 57 => (6,10,14), 58 => (6,10,14), 59 => (6,10,14), 60 => (6,10,14), 61 => (6,10,14), 62 => (6,10,14), 63 => (6,10,14), 64 => (6,10,14), 65 => (6,10,14), 66 => (6,10,14), 67 => (6,10,14), 68 => (6,10,14), 69 => (6,10,14), 70 => (5,10,14), 71 => (8,8,9), 72 => (0,0,12), 73 => (0,0,11), 74 => (1,1,12), 75 => (1,1,12), 76 => (0,0,11), 77 => (0,0,11), 78 => (0,0,11), 79 => (0,0,11), 80 => (0,0,11), 81 => (0,0,11), 82 => (0,0,11), 83 => (0,0,11), 84 => (0,0,11), 85 => (0,0,11), 86 => (0,0,11), 87 => (0,0,12), 88 => (5,5,11), 89 => (6,10,0), 90 => (9,14,0), 91 => (6,12,0), 92 => (0,9,0), 93 => (0,8,4), 94 => (4,10,11), 95 => (6,10,15), 96 => (5,10,15), 97 => (5,10,14), 98 => (5,10,15), 99 => (6,10,14), 100 => (6,10,14), 101 => (5,10,14), 102 => (5,10,14), 103 => (5,10,14), 104 => (6,10,14), 105 => (6,10,14), 106 => (6,10,15), 107 => (5,10,14), 108 => (5,10,14), 109 => (6,10,14), 110 => (6,10,14), 111 => (6,10,14), 112 => (6,10,14), 113 => (6,10,14), 114 => (6,10,14), 115 => (6,10,14), 116 => (6,10,14), 117 => (6,10,14), 118 => (6,10,14), 119 => (6,10,14), 120 => (6,10,14), 121 => (6,10,14), 122 => (6,10,15), 123 => (6,11,15), 124 => (6,11,15), 125 => (4,11,15), 126 => (9,4,7), 127 => (8,5,8), 128 => (13,0,0), 129 => (12,0,0), 130 => (12,0,0), 131 => (12,0,0), 132 => (12,0,0), 133 => (12,0,0), 134 => (7,8,11), 135 => (5,10,14), 136 => (6,10,14), 137 => (6,10,14), 138 => (6,10,14), 139 => (6,10,14), 140 => (6,10,14), 141 => (6,10,14), 142 => (6,10,14), 143 => (6,10,14), 144 => (6,10,14), 145 => (6,10,14), 146 => (6,10,14), 147 => (6,10,14), 148 => (6,10,14), 149 => (6,10,14), 150 => (6,10,14), 151 => (6,10,14), 152 => (6,10,14), 153 => (6,10,14), 154 => (6,10,14), 155 => (6,10,14), 156 => (6,10,14), 157 => (6,10,14), 158 => (6,10,14), 159 => (6,10,14)), 
			88 => (0 => (7,10,14), 1 => (7,10,14), 2 => (7,10,14), 3 => (7,10,14), 4 => (7,10,14), 5 => (7,10,14), 6 => (7,10,14), 7 => (7,10,14), 8 => (7,10,14), 9 => (7,10,14), 10 => (7,10,14), 11 => (7,10,14), 12 => (7,10,14), 13 => (7,10,14), 14 => (7,10,14), 15 => (7,10,14), 16 => (7,10,14), 17 => (7,10,14), 18 => (7,10,14), 19 => (7,10,14), 20 => (7,10,14), 21 => (7,10,14), 22 => (7,10,14), 23 => (7,10,14), 24 => (6,11,15), 25 => (11,0,0), 26 => (12,0,0), 27 => (10,1,2), 28 => (9,5,7), 29 => (10,4,6), 30 => (5,12,15), 31 => (6,11,15), 32 => (6,11,14), 33 => (6,11,14), 34 => (7,10,14), 35 => (7,10,14), 36 => (7,10,14), 37 => (7,10,14), 38 => (7,10,14), 39 => (7,10,14), 40 => (7,10,14), 41 => (7,10,14), 42 => (8,10,15), 43 => (6,10,12), 44 => (0,8,4), 45 => (0,7,0), 46 => (3,10,0), 47 => (8,13,0), 48 => (5,11,1), 49 => (7,10,15), 50 => (7,10,14), 51 => (7,10,14), 52 => (7,10,14), 53 => (7,10,14), 54 => (7,10,14), 55 => (7,10,14), 56 => (7,10,14), 57 => (7,10,14), 58 => (7,10,14), 59 => (7,10,14), 60 => (7,10,14), 61 => (7,10,14), 62 => (7,10,14), 63 => (7,10,14), 64 => (7,10,14), 65 => (8,10,15), 66 => (5,10,11), 67 => (4,9,6), 68 => (6,10,11), 69 => (6,10,15), 70 => (13,14,15), 71 => (0,0,3), 72 => (0,0,12), 73 => (0,0,11), 74 => (2,2,13), 75 => (0,0,11), 76 => (9,9,14), 77 => (8,8,14), 78 => (8,8,14), 79 => (7,7,14), 80 => (7,7,14), 81 => (6,6,14), 82 => (7,7,14), 83 => (7,7,14), 84 => (7,7,14), 85 => (6,6,14), 86 => (5,5,13), 87 => (15,15,15), 88 => (7,7,6), 89 => (5,12,3), 90 => (3,10,0), 91 => (8,13,0), 92 => (6,11,0), 93 => (7,11,0), 94 => (6,5,3), 95 => (5,5,2), 96 => (14,8,0), 97 => (15,12,8), 98 => (7,11,3), 99 => (5,11,6), 100 => (5,11,5), 101 => (8,11,15), 102 => (8,11,15), 103 => (8,11,15), 104 => (7,11,11), 105 => (5,11,6), 106 => (1,10,0), 107 => (11,10,5), 108 => (7,9,12), 109 => (6,10,14), 110 => (6,10,14), 111 => (7,10,14), 112 => (7,10,14), 113 => (7,10,14), 114 => (7,10,14), 115 => (7,10,14), 116 => (7,10,14), 117 => (7,10,14), 118 => (7,10,14), 119 => (7,10,14), 120 => (8,10,15), 121 => (6,10,11), 122 => (3,9,8), 123 => (0,7,0), 124 => (0,7,0), 125 => (7,12,0), 126 => (8,14,0), 127 => (4,11,7), 128 => (6,11,15), 129 => (6,12,15), 130 => (10,4,6), 131 => (9,5,7), 132 => (12,2,2), 133 => (12,0,0), 134 => (11,0,0), 135 => (6,11,15), 136 => (7,10,14), 137 => (7,10,14), 138 => (7,10,14), 139 => (7,10,14), 140 => (7,10,14), 141 => (7,10,14), 142 => (7,10,14), 143 => (7,10,14), 144 => (7,10,14), 145 => (7,10,14), 146 => (7,10,14), 147 => (7,10,14), 148 => (7,10,14), 149 => (7,10,14), 150 => (7,10,14), 151 => (7,10,14), 152 => (7,10,14), 153 => (7,10,14), 154 => (7,10,14), 155 => (7,10,14), 156 => (7,10,14), 157 => (7,10,14), 158 => (7,10,14), 159 => (7,10,14)), 
			89 => (0 => (7,10,14), 1 => (7,10,14), 2 => (7,10,14), 3 => (7,10,14), 4 => (7,10,14), 5 => (7,10,14), 6 => (7,10,14), 7 => (7,10,14), 8 => (7,10,14), 9 => (7,10,14), 10 => (7,10,14), 11 => (7,10,14), 12 => (7,10,14), 13 => (7,10,14), 14 => (7,10,14), 15 => (7,10,14), 16 => (7,10,14), 17 => (7,10,14), 18 => (7,10,14), 19 => (7,10,14), 20 => (7,10,14), 21 => (7,10,14), 22 => (7,10,14), 23 => (7,10,14), 24 => (7,10,14), 25 => (7,11,15), 26 => (7,12,15), 27 => (7,11,15), 28 => (7,11,14), 29 => (7,11,14), 30 => (7,10,14), 31 => (7,10,14), 32 => (7,10,14), 33 => (7,10,14), 34 => (7,10,14), 35 => (7,10,14), 36 => (7,10,14), 37 => (7,10,14), 38 => (7,10,14), 39 => (8,11,14), 40 => (8,11,15), 41 => (7,10,12), 42 => (0,8,3), 43 => (0,7,0), 44 => (0,8,1), 45 => (4,11,0), 46 => (9,13,0), 47 => (7,12,0), 48 => (11,14,0), 49 => (3,10,0), 50 => (2,8,8), 51 => (9,11,15), 52 => (8,11,15), 53 => (8,11,14), 54 => (7,10,14), 55 => (7,10,14), 56 => (7,10,14), 57 => (7,10,14), 58 => (7,10,14), 59 => (7,10,14), 60 => (8,11,14), 61 => (8,11,14), 62 => (8,11,14), 63 => (9,11,15), 64 => (3,9,7), 65 => (0,7,4), 66 => (0,8,0), 67 => (3,11,0), 68 => (5,12,0), 69 => (6,12,2), 70 => (9,12,12), 71 => (0,0,4), 72 => (0,0,12), 73 => (1,1,12), 74 => (1,1,12), 75 => (0,0,12), 76 => (0,0,3), 77 => (0,0,4), 78 => (0,0,4), 79 => (0,0,4), 80 => (0,0,4), 81 => (0,0,4), 82 => (0,0,4), 83 => (0,0,4), 84 => (0,0,4), 85 => (0,0,4), 86 => (0,0,4), 87 => (0,0,4), 88 => (0,0,1), 89 => (9,13,9), 90 => (2,9,0), 91 => (2,9,1), 92 => (2,10,1), 93 => (0,8,1), 94 => (7,8,1), 95 => (7,7,3), 96 => (10,7,3), 97 => (13,11,6), 98 => (15,12,9), 99 => (9,9,3), 100 => (11,7,3), 101 => (9,5,1), 102 => (9,11,2), 103 => (5,11,3), 104 => (1,10,0), 105 => (11,9,3), 106 => (15,12,9), 107 => (14,12,8), 108 => (14,11,6), 109 => (14,11,7), 110 => (8,10,12), 111 => (7,11,14), 112 => (7,10,14), 113 => (7,10,14), 114 => (7,10,14), 115 => (7,10,14), 116 => (8,11,14), 117 => (9,11,15), 118 => (7,10,11), 119 => (4,9,8), 120 => (0,8,4), 121 => (0,7,0), 122 => (0,7,1), 123 => (0,8,1), 124 => (1,9,0), 125 => (1,9,0), 126 => (7,12,0), 127 => (9,14,0), 128 => (9,14,0), 129 => (6,11,7), 130 => (7,11,15), 131 => (7,11,15), 132 => (7,11,15), 133 => (7,12,15), 134 => (7,11,15), 135 => (7,10,14), 136 => (7,10,14), 137 => (7,10,14), 138 => (7,10,14), 139 => (7,10,14), 140 => (7,10,14), 141 => (7,10,14), 142 => (7,10,14), 143 => (7,10,14), 144 => (7,10,14), 145 => (7,10,14), 146 => (7,10,14), 147 => (7,10,14), 148 => (7,10,14), 149 => (7,10,14), 150 => (7,10,14), 151 => (7,10,14), 152 => (7,10,14), 153 => (7,10,14), 154 => (7,10,14), 155 => (7,10,14), 156 => (7,10,14), 157 => (7,10,14), 158 => (7,10,14), 159 => (7,10,14)), 
			90 => (0 => (10,12,14), 1 => (10,12,14), 2 => (10,12,14), 3 => (10,12,14), 4 => (10,12,14), 5 => (10,12,14), 6 => (10,12,14), 7 => (10,12,14), 8 => (10,12,14), 9 => (10,12,14), 10 => (10,12,14), 11 => (10,12,14), 12 => (10,12,14), 13 => (10,12,14), 14 => (10,12,14), 15 => (10,12,14), 16 => (10,12,14), 17 => (10,12,14), 18 => (10,12,14), 19 => (10,12,14), 20 => (10,12,14), 21 => (10,12,14), 22 => (10,12,14), 23 => (10,12,14), 24 => (10,12,14), 25 => (10,12,14), 26 => (10,12,14), 27 => (10,12,14), 28 => (10,12,14), 29 => (10,12,14), 30 => (10,12,14), 31 => (10,12,14), 32 => (10,12,14), 33 => (10,12,14), 34 => (11,12,15), 35 => (11,12,15), 36 => (11,12,15), 37 => (10,12,14), 38 => (11,12,15), 39 => (8,11,11), 40 => (5,10,8), 41 => (0,8,0), 42 => (0,8,1), 43 => (1,9,0), 44 => (0,7,1), 45 => (4,11,0), 46 => (5,11,0), 47 => (9,13,0), 48 => (9,13,0), 49 => (10,14,0), 50 => (7,12,0), 51 => (3,10,0), 52 => (0,8,0), 53 => (5,10,7), 54 => (11,12,15), 55 => (10,12,15), 56 => (10,12,14), 57 => (10,12,14), 58 => (10,12,15), 59 => (11,12,15), 60 => (4,9,7), 61 => (5,10,8), 62 => (5,10,8), 63 => (0,7,0), 64 => (0,7,1), 65 => (0,9,0), 66 => (4,11,0), 67 => (7,12,0), 68 => (9,13,0), 69 => (6,12,0), 70 => (11,15,7), 71 => (0,0,5), 72 => (0,0,12), 73 => (2,2,13), 74 => (0,0,11), 75 => (0,0,12), 76 => (0,0,12), 77 => (0,0,12), 78 => (0,0,12), 79 => (0,0,12), 80 => (0,0,12), 81 => (0,0,12), 82 => (0,0,12), 83 => (0,0,12), 84 => (0,0,12), 85 => (0,0,12), 86 => (0,0,12), 87 => (0,0,13), 88 => (0,0,5), 89 => (9,14,7), 90 => (0,7,1), 91 => (0,7,2), 92 => (10,7,0), 93 => (11,11,3), 94 => (4,13,0), 95 => (2,9,0), 96 => (8,5,2), 97 => (13,8,0), 98 => (8,11,1), 99 => (11,10,1), 100 => (10,6,1), 101 => (5,6,3), 102 => (5,12,0), 103 => (7,13,0), 104 => (13,13,4), 105 => (11,11,0), 106 => (10,6,1), 107 => (14,10,7), 108 => (14,11,8), 109 => (14,11,7), 110 => (14,11,7), 111 => (15,11,8), 112 => (10,12,7), 113 => (11,13,11), 114 => (15,15,15), 115 => (12,13,11), 116 => (7,12,7), 117 => (0,7,0), 118 => (0,7,0), 119 => (0,7,1), 120 => (0,7,1), 121 => (0,7,2), 122 => (0,8,1), 123 => (2,10,0), 124 => (0,7,2), 125 => (0,8,1), 126 => (3,10,0), 127 => (6,12,0), 128 => (10,14,0), 129 => (7,12,0), 130 => (7,13,0), 131 => (10,13,7), 132 => (10,11,15), 133 => (10,12,14), 134 => (10,12,14), 135 => (10,12,14), 136 => (10,12,14), 137 => (10,12,14), 138 => (10,12,14), 139 => (10,12,14), 140 => (10,12,14), 141 => (10,12,14), 142 => (10,12,14), 143 => (10,12,14), 144 => (10,12,14), 145 => (10,12,14), 146 => (10,12,14), 147 => (10,12,14), 148 => (10,12,14), 149 => (10,12,14), 150 => (10,12,14), 151 => (10,12,14), 152 => (10,12,14), 153 => (10,12,14), 154 => (10,12,14), 155 => (10,12,14), 156 => (10,12,14), 157 => (10,12,14), 158 => (10,12,14), 159 => (10,12,14)), 
			91 => (0 => (9,11,14), 1 => (9,11,14), 2 => (9,11,14), 3 => (9,11,14), 4 => (9,11,14), 5 => (9,11,14), 6 => (9,11,14), 7 => (9,11,14), 8 => (9,11,14), 9 => (9,11,14), 10 => (9,11,14), 11 => (9,11,14), 12 => (9,11,14), 13 => (9,11,14), 14 => (9,11,14), 15 => (9,11,14), 16 => (9,11,14), 17 => (9,11,14), 18 => (9,11,14), 19 => (9,11,14), 20 => (9,11,14), 21 => (10,12,14), 22 => (9,11,14), 23 => (9,11,14), 24 => (9,11,14), 25 => (9,11,14), 26 => (9,11,14), 27 => (9,11,14), 28 => (9,11,14), 29 => (9,11,14), 30 => (9,11,14), 31 => (10,12,14), 32 => (11,12,15), 33 => (4,9,7), 34 => (1,8,4), 35 => (0,7,0), 36 => (1,8,4), 37 => (5,10,9), 38 => (0,7,0), 39 => (0,8,0), 40 => (0,9,0), 41 => (0,7,2), 42 => (1,9,0), 43 => (1,9,0), 44 => (3,10,1), 45 => (4,11,0), 46 => (4,11,0), 47 => (5,11,0), 48 => (6,12,0), 49 => (4,11,0), 50 => (11,14,0), 51 => (9,13,0), 52 => (8,13,0), 53 => (5,12,0), 54 => (2,10,0), 55 => (5,11,2), 56 => (6,10,8), 57 => (4,9,8), 58 => (5,11,3), 59 => (0,8,0), 60 => (0,9,0), 61 => (0,8,0), 62 => (0,8,0), 63 => (1,10,0), 64 => (2,10,0), 65 => (5,11,0), 66 => (5,11,0), 67 => (9,13,0), 68 => (10,14,0), 69 => (6,12,0), 70 => (10,12,8), 71 => (0,0,5), 72 => (1,1,13), 73 => (1,1,12), 74 => (0,0,11), 75 => (0,0,12), 76 => (0,0,12), 77 => (0,0,12), 78 => (0,0,12), 79 => (0,0,12), 80 => (0,0,12), 81 => (0,0,12), 82 => (0,0,12), 83 => (0,0,12), 84 => (0,0,12), 85 => (0,0,12), 86 => (0,0,12), 87 => (0,0,12), 88 => (0,0,5), 89 => (11,11,8), 90 => (3,9,0), 91 => (7,8,0), 92 => (13,8,0), 93 => (15,10,8), 94 => (12,10,4), 95 => (15,10,6), 96 => (15,11,9), 97 => (12,11,6), 98 => (10,11,3), 99 => (9,10,0), 100 => (9,6,5), 101 => (7,10,2), 102 => (7,11,4), 103 => (11,10,5), 104 => (11,11,7), 105 => (3,7,4), 106 => (13,9,5), 107 => (10,6,0), 108 => (14,9,5), 109 => (12,7,0), 110 => (14,9,5), 111 => (12,10,6), 112 => (15,11,6), 113 => (6,8,0), 114 => (0,8,0), 115 => (0,8,0), 116 => (9,4,4), 117 => (1,7,2), 118 => (0,7,2), 119 => (0,7,2), 120 => (0,8,2), 121 => (0,7,2), 122 => (0,8,0), 123 => (5,11,0), 124 => (0,7,2), 125 => (1,9,0), 126 => (4,11,0), 127 => (7,12,0), 128 => (11,14,0), 129 => (11,14,0), 130 => (9,13,0), 131 => (10,14,0), 132 => (10,14,0), 133 => (10,13,7), 134 => (10,12,15), 135 => (10,11,14), 136 => (9,11,14), 137 => (9,11,14), 138 => (9,11,14), 139 => (9,11,14), 140 => (9,11,14), 141 => (9,11,14), 142 => (9,11,14), 143 => (9,11,14), 144 => (9,11,14), 145 => (9,11,14), 146 => (9,11,14), 147 => (9,11,14), 148 => (9,11,14), 149 => (9,11,14), 150 => (9,11,14), 151 => (9,11,14), 152 => (9,11,14), 153 => (9,11,14), 154 => (9,11,14), 155 => (9,11,14), 156 => (9,11,14), 157 => (9,11,14), 158 => (9,11,14), 159 => (9,11,14)), 
			92 => (0 => (12,13,14), 1 => (12,13,14), 2 => (12,13,14), 3 => (12,13,14), 4 => (12,13,14), 5 => (12,13,14), 6 => (12,13,14), 7 => (12,13,14), 8 => (12,13,14), 9 => (12,13,14), 10 => (12,13,14), 11 => (12,13,14), 12 => (12,13,14), 13 => (12,13,14), 14 => (12,13,14), 15 => (12,13,14), 16 => (12,13,14), 17 => (12,13,14), 18 => (12,13,14), 19 => (12,13,14), 20 => (14,13,15), 21 => (4,9,7), 22 => (12,14,6), 23 => (11,13,11), 24 => (13,13,15), 25 => (13,13,15), 26 => (13,13,14), 27 => (13,13,14), 28 => (13,13,14), 29 => (13,13,15), 30 => (14,14,15), 31 => (6,10,8), 32 => (0,7,0), 33 => (0,7,1), 34 => (0,7,1), 35 => (0,7,2), 36 => (1,9,0), 37 => (0,7,1), 38 => (0,9,0), 39 => (0,8,0), 40 => (0,8,1), 41 => (0,7,2), 42 => (0,7,2), 43 => (0,8,1), 44 => (0,7,1), 45 => (1,9,0), 46 => (6,12,0), 47 => (8,13,0), 48 => (8,13,0), 49 => (6,12,0), 50 => (9,13,0), 51 => (10,14,0), 52 => (11,14,0), 53 => (7,12,0), 54 => (6,12,0), 55 => (4,11,0), 56 => (4,11,0), 57 => (4,12,0), 58 => (3,11,0), 59 => (0,9,0), 60 => (3,11,0), 61 => (5,11,0), 62 => (5,11,0), 63 => (6,12,0), 64 => (8,13,0), 65 => (4,11,0), 66 => (7,12,0), 67 => (10,14,0), 68 => (9,13,0), 69 => (2,10,0), 70 => (8,12,7), 71 => (0,0,4), 72 => (0,0,13), 73 => (0,0,11), 74 => (0,0,11), 75 => (0,0,11), 76 => (0,0,11), 77 => (0,0,11), 78 => (0,0,11), 79 => (0,0,11), 80 => (0,0,11), 81 => (0,0,11), 82 => (0,0,11), 83 => (0,0,11), 84 => (0,0,11), 85 => (0,0,11), 86 => (0,0,11), 87 => (0,0,12), 88 => (0,0,4), 89 => (9,10,7), 90 => (5,7,0), 91 => (2,8,0), 92 => (14,9,3), 93 => (12,9,3), 94 => (13,10,5), 95 => (13,7,1), 96 => (12,11,7), 97 => (9,10,2), 98 => (6,11,0), 99 => (7,12,1), 100 => (14,10,10), 101 => (15,10,6), 102 => (9,9,4), 103 => (10,10,4), 104 => (0,9,5), 105 => (5,7,3), 106 => (5,9,2), 107 => (14,10,7), 108 => (4,8,2), 109 => (6,8,0), 110 => (10,8,0), 111 => (9,6,5), 112 => (9,5,4), 113 => (11,11,6), 114 => (13,6,4), 115 => (7,11,0), 116 => (5,13,0), 117 => (9,8,2), 118 => (1,9,1), 119 => (3,10,0), 120 => (0,7,2), 121 => (0,7,2), 122 => (5,11,0), 123 => (7,12,0), 124 => (2,9,1), 125 => (0,7,1), 126 => (2,9,1), 127 => (8,13,0), 128 => (4,11,0), 129 => (3,10,0), 130 => (6,12,0), 131 => (7,12,0), 132 => (7,12,0), 133 => (8,13,0), 134 => (1,10,0), 135 => (11,12,12), 136 => (13,13,15), 137 => (12,13,14), 138 => (12,13,14), 139 => (12,13,14), 140 => (12,13,14), 141 => (12,13,14), 142 => (12,13,14), 143 => (12,13,14), 144 => (12,13,14), 145 => (12,13,14), 146 => (12,13,14), 147 => (12,13,14), 148 => (12,13,14), 149 => (12,13,14), 150 => (12,13,14), 151 => (12,13,14), 152 => (12,13,14), 153 => (12,13,14), 154 => (12,13,14), 155 => (12,13,14), 156 => (12,13,14), 157 => (12,13,14), 158 => (12,13,14), 159 => (12,13,14)), 
			93 => (0 => (13,13,14), 1 => (13,13,14), 2 => (13,13,14), 3 => (13,13,14), 4 => (13,13,14), 5 => (13,13,14), 6 => (13,13,14), 7 => (13,13,14), 8 => (13,13,14), 9 => (13,13,14), 10 => (13,13,14), 11 => (13,13,14), 12 => (13,13,14), 13 => (13,13,14), 14 => (13,13,14), 15 => (13,13,14), 16 => (13,13,14), 17 => (14,14,15), 18 => (15,14,15), 19 => (8,12,7), 20 => (0,8,0), 21 => (6,12,0), 22 => (6,12,0), 23 => (10,14,0), 24 => (3,10,0), 25 => (3,10,0), 26 => (5,9,9), 27 => (5,10,8), 28 => (6,10,8), 29 => (3,9,3), 30 => (0,7,0), 31 => (0,7,1), 32 => (0,8,2), 33 => (0,7,2), 34 => (0,8,1), 35 => (1,10,0), 36 => (0,8,1), 37 => (0,7,2), 38 => (4,11,0), 39 => (7,12,0), 40 => (0,7,2), 41 => (0,8,1), 42 => (0,7,2), 43 => (0,8,1), 44 => (8,13,0), 45 => (4,11,0), 46 => (8,13,0), 47 => (9,13,0), 48 => (11,14,0), 49 => (5,11,0), 50 => (8,13,0), 51 => (8,13,0), 52 => (5,12,0), 53 => (2,10,0), 54 => (4,9,0), 55 => (7,9,0), 56 => (10,8,0), 57 => (10,5,1), 58 => (10,8,0), 59 => (10,9,5), 60 => (9,9,0), 61 => (7,11,0), 62 => (5,10,0), 63 => (7,13,0), 64 => (5,12,0), 65 => (5,12,0), 66 => (6,12,0), 67 => (7,13,0), 68 => (5,12,0), 69 => (9,14,0), 70 => (13,15,8), 71 => (5,5,11), 72 => (6,6,15), 73 => (6,6,14), 74 => (6,6,14), 75 => (6,6,14), 76 => (6,6,14), 77 => (6,6,14), 78 => (6,6,14), 79 => (6,6,14), 80 => (6,6,14), 81 => (6,6,14), 82 => (6,6,14), 83 => (6,6,14), 84 => (6,6,14), 85 => (6,6,14), 86 => (6,6,14), 87 => (6,6,15), 88 => (5,5,11), 89 => (13,12,13), 90 => (14,9,2), 91 => (5,10,7), 92 => (4,10,8), 93 => (13,10,6), 94 => (14,11,7), 95 => (11,13,8), 96 => (6,13,3), 97 => (9,10,0), 98 => (14,8,3), 99 => (9,10,0), 100 => (5,10,1), 101 => (5,10,1), 102 => (11,10,7), 103 => (10,8,3), 104 => (10,9,3), 105 => (9,8,0), 106 => (9,5,3), 107 => (6,7,2), 108 => (7,10,3), 109 => (5,13,0), 110 => (2,11,0), 111 => (1,10,0), 112 => (3,11,0), 113 => (3,10,0), 114 => (0,9,1), 115 => (5,8,0), 116 => (2,10,1), 117 => (0,8,1), 118 => (0,6,2), 119 => (8,13,0), 120 => (6,12,0), 121 => (2,10,0), 122 => (3,10,0), 123 => (6,12,0), 124 => (7,12,0), 125 => (2,10,0), 126 => (1,10,0), 127 => (0,9,0), 128 => (0,8,1), 129 => (0,9,0), 130 => (0,8,1), 131 => (0,9,0), 132 => (2,10,0), 133 => (5,11,0), 134 => (5,11,0), 135 => (4,11,0), 136 => (5,11,2), 137 => (6,11,7), 138 => (10,12,11), 139 => (14,13,15), 140 => (14,13,15), 141 => (13,13,14), 142 => (13,13,14), 143 => (13,13,14), 144 => (13,13,14), 145 => (13,13,14), 146 => (13,13,14), 147 => (13,13,14), 148 => (13,13,14), 149 => (13,13,14), 150 => (13,13,14), 151 => (13,13,14), 152 => (13,13,14), 153 => (13,13,14), 154 => (13,13,14), 155 => (13,13,14), 156 => (13,13,14), 157 => (13,13,14), 158 => (13,13,14), 159 => (13,13,14)), 
			94 => (0 => (14,14,14), 1 => (14,14,14), 2 => (14,14,14), 3 => (14,14,14), 4 => (14,14,14), 5 => (14,14,14), 6 => (14,14,14), 7 => (14,14,14), 8 => (14,14,14), 9 => (14,14,14), 10 => (14,14,14), 11 => (14,14,14), 12 => (14,14,14), 13 => (15,14,14), 14 => (15,14,15), 15 => (15,15,15), 16 => (6,10,7), 17 => (2,9,4), 18 => (0,8,0), 19 => (5,12,0), 20 => (4,10,1), 21 => (0,9,0), 22 => (2,10,0), 23 => (4,11,0), 24 => (11,14,0), 25 => (10,14,0), 26 => (10,14,0), 27 => (5,11,0), 28 => (0,7,0), 29 => (1,9,0), 30 => (0,8,1), 31 => (0,8,1), 32 => (0,7,2), 33 => (1,9,0), 34 => (0,8,0), 35 => (0,8,1), 36 => (2,9,1), 37 => (8,13,0), 38 => (10,14,0), 39 => (3,10,0), 40 => (1,9,0), 41 => (0,8,0), 42 => (8,13,0), 43 => (6,12,0), 44 => (8,13,0), 45 => (8,13,0), 46 => (6,12,0), 47 => (5,12,0), 48 => (1,9,0), 49 => (3,11,0), 50 => (1,10,0), 51 => (4,6,2), 52 => (7,9,3), 53 => (10,9,2), 54 => (15,12,10), 55 => (14,11,6), 56 => (14,13,11), 57 => (14,13,10), 58 => (11,7,2), 59 => (14,12,8), 60 => (13,11,7), 61 => (14,11,8), 62 => (12,9,6), 63 => (8,4,2), 64 => (6,6,2), 65 => (6,11,0), 66 => (11,8,2), 67 => (10,10,0), 68 => (10,11,0), 69 => (14,8,1), 70 => (0,5,0), 71 => (0,0,0), 72 => (0,0,0), 73 => (0,0,0), 74 => (0,0,0), 75 => (0,0,0), 76 => (0,0,0), 77 => (0,0,0), 78 => (0,0,0), 79 => (0,0,0), 80 => (0,0,0), 81 => (0,0,0), 82 => (0,0,0), 83 => (0,0,0), 84 => (0,0,0), 85 => (0,0,0), 86 => (0,0,0), 87 => (0,0,0), 88 => (0,0,0), 89 => (7,8,4), 90 => (10,8,3), 91 => (15,11,7), 92 => (15,14,15), 93 => (14,12,10), 94 => (13,11,7), 95 => (15,10,7), 96 => (9,8,0), 97 => (9,5,1), 98 => (15,13,11), 99 => (11,11,5), 100 => (6,8,0), 101 => (0,10,0), 102 => (0,10,0), 103 => (6,8,0), 104 => (15,8,3), 105 => (11,7,0), 106 => (8,5,3), 107 => (11,7,0), 108 => (10,6,1), 109 => (7,6,4), 110 => (6,11,0), 111 => (1,9,1), 112 => (2,10,0), 113 => (0,9,0), 114 => (0,9,0), 115 => (0,8,1), 116 => (0,9,1), 117 => (7,13,0), 118 => (2,10,0), 119 => (4,11,0), 120 => (0,8,1), 121 => (1,9,0), 122 => (6,12,0), 123 => (2,9,1), 124 => (4,11,0), 125 => (4,11,0), 126 => (0,9,0), 127 => (0,6,2), 128 => (4,7,1), 129 => (3,6,3), 130 => (0,8,2), 131 => (0,7,2), 132 => (0,8,1), 133 => (1,10,0), 134 => (4,9,0), 135 => (1,7,1), 136 => (0,9,0), 137 => (3,11,0), 138 => (2,11,0), 139 => (3,11,0), 140 => (3,11,1), 141 => (15,14,15), 142 => (15,14,15), 143 => (14,14,14), 144 => (14,14,14), 145 => (14,14,14), 146 => (14,14,14), 147 => (14,14,14), 148 => (14,14,14), 149 => (14,14,14), 150 => (14,14,14), 151 => (14,14,14), 152 => (14,14,14), 153 => (14,14,14), 154 => (14,14,14), 155 => (14,14,14), 156 => (14,14,14), 157 => (14,14,14), 158 => (14,14,14), 159 => (14,14,14)), 
			95 => (0 => (15,14,14), 1 => (15,15,14), 2 => (15,14,14), 3 => (15,14,14), 4 => (15,14,14), 5 => (15,15,14), 6 => (15,14,14), 7 => (15,14,14), 8 => (15,14,14), 9 => (15,15,14), 10 => (15,14,14), 11 => (15,15,14), 12 => (10,13,10), 13 => (6,11,6), 14 => (2,9,2), 15 => (0,7,0), 16 => (0,7,0), 17 => (0,8,0), 18 => (0,7,0), 19 => (0,9,0), 20 => (0,7,0), 21 => (0,8,0), 22 => (0,8,0), 23 => (0,8,0), 24 => (0,7,0), 25 => (1,10,0), 26 => (0,9,0), 27 => (0,8,0), 28 => (0,9,0), 29 => (1,9,0), 30 => (1,10,0), 31 => (1,10,0), 32 => (2,10,0), 33 => (1,10,0), 34 => (8,11,0), 35 => (12,11,2), 36 => (4,12,0), 37 => (4,12,0), 38 => (9,11,0), 39 => (6,10,0), 40 => (7,11,0), 41 => (12,12,2), 42 => (8,9,2), 43 => (8,10,1), 44 => (8,10,2), 45 => (8,9,2), 46 => (8,10,2), 47 => (8,9,0), 48 => (3,9,0), 49 => (9,10,2), 50 => (6,8,2), 51 => (0,10,0), 52 => (15,11,6), 53 => (15,12,8), 54 => (10,11,4), 55 => (15,9,5), 56 => (10,10,4), 57 => (14,15,15), 58 => (15,12,8), 59 => (14,12,9), 60 => (14,13,12), 61 => (15,14,13), 62 => (13,11,7), 63 => (13,9,2), 64 => (14,13,10), 65 => (15,12,10), 66 => (15,13,9), 67 => (15,12,7), 68 => (10,12,8), 69 => (9,10,5), 70 => (10,7,0), 71 => (0,6,0), 72 => (2,3,0), 73 => (0,5,0), 74 => (0,4,0), 75 => (0,3,0), 76 => (0,3,0), 77 => (0,3,0), 78 => (0,3,0), 79 => (0,5,0), 80 => (3,6,0), 81 => (2,6,0), 82 => (5,5,1), 83 => (4,5,0), 84 => (6,3,0), 85 => (6,4,0), 86 => (6,3,0), 87 => (1,3,0), 88 => (4,7,0), 89 => (4,12,0), 90 => (0,10,0), 91 => (4,8,2), 92 => (12,6,0), 93 => (15,12,6), 94 => (11,8,0), 95 => (10,6,0), 96 => (7,5,3), 97 => (9,6,1), 98 => (14,11,6), 99 => (15,12,8), 100 => (15,12,9), 101 => (15,11,7), 102 => (14,8,0), 103 => (11,11,3), 104 => (7,12,3), 105 => (5,9,1), 106 => (15,11,3), 107 => (10,7,3), 108 => (11,8,3), 109 => (12,7,0), 110 => (10,8,0), 111 => (10,10,0), 112 => (11,8,3), 113 => (14,10,1), 114 => (7,9,2), 115 => (4,9,0), 116 => (8,9,0), 117 => (8,9,0), 118 => (4,9,1), 119 => (0,7,0), 120 => (0,8,0), 121 => (0,9,0), 122 => (0,8,0), 123 => (0,8,0), 124 => (1,7,1), 125 => (3,6,1), 126 => (8,7,3), 127 => (13,8,4), 128 => (15,10,3), 129 => (15,9,1), 130 => (13,7,0), 131 => (8,6,1), 132 => (1,7,1), 133 => (3,8,2), 134 => (11,9,2), 135 => (14,8,3), 136 => (8,7,3), 137 => (7,6,0), 138 => (13,7,5), 139 => (11,6,0), 140 => (9,7,0), 141 => (4,10,0), 142 => (0,9,0), 143 => (8,12,5), 144 => (11,13,9), 145 => (15,15,14), 146 => (15,14,14), 147 => (15,14,14), 148 => (15,14,14), 149 => (15,15,14), 150 => (15,14,14), 151 => (15,14,14), 152 => (15,14,14), 153 => (15,15,14), 154 => (15,14,14), 155 => (15,14,14), 156 => (15,14,14), 157 => (15,15,14), 158 => (15,14,14), 159 => (15,14,14)), 
			96 => (0 => (3,6,14), 1 => (2,5,14), 2 => (4,7,14), 3 => (3,5,14), 4 => (3,5,14), 5 => (2,5,14), 6 => (5,7,14), 7 => (3,6,14), 8 => (3,6,14), 9 => (2,5,14), 10 => (5,8,14), 11 => (3,6,14), 12 => (3,6,14), 13 => (3,5,14), 14 => (5,8,15), 15 => (4,6,15), 16 => (4,6,15), 17 => (3,5,15), 18 => (6,8,15), 19 => (5,7,15), 20 => (5,6,15), 21 => (4,6,15), 22 => (3,5,15), 23 => (6,8,15), 24 => (5,7,15), 25 => (4,6,15), 26 => (3,5,15), 27 => (7,8,15), 28 => (4,6,15), 29 => (3,5,15), 30 => (6,8,15), 31 => (4,6,15), 32 => (4,6,15), 33 => (3,5,15), 34 => (6,8,15), 35 => (4,6,15), 36 => (4,6,15), 37 => (3,5,15), 38 => (5,7,15), 39 => (3,6,15), 40 => (3,6,15), 41 => (2,5,15), 42 => (5,8,15), 43 => (4,7,15), 44 => (3,6,15), 45 => (6,8,15), 46 => (4,5,15), 47 => (4,6,15), 48 => (4,6,15), 49 => (1,3,15), 50 => (14,14,15), 51 => (5,5,15), 52 => (10,9,12), 53 => (8,1,2), 54 => (9,1,2), 55 => (11,9,12), 56 => (8,9,15), 57 => (13,13,14), 58 => (4,7,14), 59 => (7,10,14), 60 => (15,15,14), 61 => (3,5,14), 62 => (13,14,10), 63 => (9,11,7), 64 => (7,7,6), 65 => (6,8,15), 66 => (8,11,14), 67 => (2,5,14), 68 => (2,4,14), 69 => (9,11,15), 70 => (15,15,7), 71 => (13,13,8), 72 => (12,13,8), 73 => (5,6,14), 74 => (12,12,8), 75 => (9,10,7), 76 => (10,12,15), 77 => (8,9,15), 78 => (7,9,15), 79 => (10,11,7), 80 => (6,6,7), 81 => (6,9,15), 82 => (13,14,7), 83 => (5,6,8), 84 => (10,12,8), 85 => (5,7,8), 86 => (9,11,8), 87 => (12,14,8), 88 => (11,12,8), 89 => (6,6,7), 90 => (10,11,8), 91 => (12,14,8), 92 => (9,11,8), 93 => (0,2,12), 94 => (5,8,15), 95 => (4,7,15), 96 => (4,7,15), 97 => (2,6,15), 98 => (4,7,14), 99 => (3,6,14), 100 => (3,6,14), 101 => (2,5,14), 102 => (5,8,15), 103 => (4,6,15), 104 => (4,6,15), 105 => (3,5,15), 106 => (2,5,15), 107 => (5,8,15), 108 => (4,7,15), 109 => (3,6,15), 110 => (2,5,15), 111 => (6,8,15), 112 => (3,6,15), 113 => (2,5,15), 114 => (5,8,15), 115 => (4,6,15), 116 => (3,6,15), 117 => (2,5,15), 118 => (6,8,15), 119 => (5,7,15), 120 => (4,6,15), 121 => (3,5,15), 122 => (6,8,15), 123 => (4,6,15), 124 => (4,6,15), 125 => (3,5,15), 126 => (5,8,15), 127 => (4,7,15), 128 => (3,6,15), 129 => (2,5,15), 130 => (5,8,15), 131 => (3,6,15), 132 => (4,6,15), 133 => (3,5,15), 134 => (5,8,15), 135 => (3,7,15), 136 => (4,6,15), 137 => (3,5,15), 138 => (5,8,15), 139 => (3,6,15), 140 => (3,6,15), 141 => (3,5,15), 142 => (6,8,15), 143 => (4,6,14), 144 => (3,6,14), 145 => (2,5,14), 146 => (4,7,14), 147 => (3,5,14), 148 => (3,5,14), 149 => (2,5,14), 150 => (5,7,14), 151 => (3,6,14), 152 => (3,6,14), 153 => (2,5,14), 154 => (4,7,14), 155 => (3,5,14), 156 => (3,5,14), 157 => (2,5,14), 158 => (5,7,14), 159 => (3,6,14)), 
			97 => (0 => (0,1,14), 1 => (1,3,14), 2 => (1,3,14), 3 => (0,2,14), 4 => (2,4,14), 5 => (1,3,14), 6 => (3,6,14), 7 => (1,3,14), 8 => (0,1,14), 9 => (0,2,14), 10 => (2,4,14), 11 => (1,3,14), 12 => (0,1,14), 13 => (1,3,14), 14 => (1,3,14), 15 => (0,2,14), 16 => (2,4,14), 17 => (1,3,14), 18 => (3,6,14), 19 => (1,3,14), 20 => (0,1,14), 21 => (1,3,14), 22 => (3,6,14), 23 => (0,2,14), 24 => (2,4,14), 25 => (0,2,14), 26 => (1,3,14), 27 => (1,3,14), 28 => (0,1,14), 29 => (1,3,14), 30 => (1,3,14), 31 => (0,2,14), 32 => (2,4,14), 33 => (1,3,14), 34 => (3,6,14), 35 => (1,3,14), 36 => (0,1,14), 37 => (1,3,14), 38 => (1,3,14), 39 => (0,2,14), 40 => (2,4,14), 41 => (1,3,14), 42 => (3,6,14), 43 => (1,3,14), 44 => (0,1,14), 45 => (0,2,14), 46 => (4,6,14), 47 => (4,6,14), 48 => (4,7,14), 49 => (6,10,14), 50 => (5,5,14), 51 => (15,15,15), 52 => (8,0,0), 53 => (11,10,4), 54 => (11,10,4), 55 => (8,0,0), 56 => (15,15,15), 57 => (10,12,14), 58 => (1,3,14), 59 => (9,11,14), 60 => (5,8,14), 61 => (8,10,14), 62 => (6,8,15), 63 => (15,15,0), 64 => (6,5,0), 65 => (7,9,15), 66 => (4,6,14), 67 => (6,8,14), 68 => (5,7,14), 69 => (7,8,15), 70 => (15,15,0), 71 => (4,4,0), 72 => (15,15,0), 73 => (6,5,0), 74 => (15,15,0), 75 => (6,5,0), 76 => (4,7,15), 77 => (4,6,14), 78 => (4,6,11), 79 => (11,11,0), 80 => (11,9,0), 81 => (0,0,13), 82 => (13,13,1), 83 => (4,4,0), 84 => (15,15,0), 85 => (1,1,2), 86 => (15,15,0), 87 => (11,11,0), 88 => (2,2,0), 89 => (0,0,7), 90 => (15,15,0), 91 => (4,4,0), 92 => (15,15,0), 93 => (7,6,0), 94 => (2,5,15), 95 => (1,3,14), 96 => (0,1,14), 97 => (1,3,14), 98 => (1,3,14), 99 => (0,2,14), 100 => (2,4,14), 101 => (1,3,14), 102 => (3,6,14), 103 => (1,3,14), 104 => (0,1,14), 105 => (1,3,14), 106 => (3,6,14), 107 => (0,2,14), 108 => (2,4,14), 109 => (0,2,14), 110 => (1,3,14), 111 => (1,3,14), 112 => (0,1,14), 113 => (1,3,14), 114 => (1,3,14), 115 => (0,2,14), 116 => (2,4,14), 117 => (1,3,14), 118 => (3,6,14), 119 => (1,3,14), 120 => (0,1,14), 121 => (1,3,14), 122 => (1,3,14), 123 => (0,2,14), 124 => (2,4,14), 125 => (1,3,14), 126 => (3,6,14), 127 => (1,3,14), 128 => (0,1,14), 129 => (1,3,14), 130 => (1,3,14), 131 => (0,2,14), 132 => (2,4,14), 133 => (1,3,14), 134 => (3,6,14), 135 => (1,3,14), 136 => (0,1,14), 137 => (1,3,14), 138 => (1,3,14), 139 => (0,2,14), 140 => (2,4,14), 141 => (1,3,14), 142 => (3,6,14), 143 => (1,3,14), 144 => (0,1,14), 145 => (1,3,14), 146 => (1,3,14), 147 => (0,2,14), 148 => (2,4,14), 149 => (1,3,14), 150 => (3,6,14), 151 => (1,3,14), 152 => (0,1,14), 153 => (1,3,14), 154 => (1,3,14), 155 => (0,2,14), 156 => (2,4,14), 157 => (1,3,14), 158 => (3,6,14), 159 => (1,2,14)), 
			98 => (0 => (0,2,14), 1 => (0,1,14), 2 => (0,1,14), 3 => (1,3,14), 4 => (0,1,14), 5 => (0,1,14), 6 => (0,1,14), 7 => (1,3,14), 8 => (0,1,14), 9 => (0,1,14), 10 => (0,1,14), 11 => (0,1,14), 12 => (0,2,14), 13 => (0,1,14), 14 => (0,1,14), 15 => (1,3,14), 16 => (0,1,14), 17 => (0,1,14), 18 => (0,1,14), 19 => (1,3,14), 20 => (0,1,14), 21 => (1,3,14), 22 => (0,1,14), 23 => (0,1,14), 24 => (0,1,14), 25 => (0,1,14), 26 => (1,3,14), 27 => (0,1,14), 28 => (0,2,14), 29 => (0,1,14), 30 => (0,1,14), 31 => (1,3,14), 32 => (0,1,14), 33 => (0,1,14), 34 => (0,1,14), 35 => (1,3,14), 36 => (0,1,14), 37 => (0,1,14), 38 => (0,1,14), 39 => (1,3,14), 40 => (0,1,14), 41 => (0,1,14), 42 => (0,1,14), 43 => (1,3,14), 44 => (0,2,14), 45 => (1,3,14), 46 => (4,6,14), 47 => (0,1,14), 48 => (5,6,14), 49 => (3,5,14), 50 => (6,7,14), 51 => (14,14,15), 52 => (7,0,0), 53 => (8,6,0), 54 => (8,6,0), 55 => (7,0,0), 56 => (14,14,15), 57 => (0,0,14), 58 => (10,13,14), 59 => (8,9,14), 60 => (5,7,14), 61 => (11,13,14), 62 => (6,8,15), 63 => (15,15,0), 64 => (6,6,0), 65 => (5,7,15), 66 => (8,10,14), 67 => (1,3,14), 68 => (1,3,14), 69 => (0,2,15), 70 => (15,15,0), 71 => (11,11,0), 72 => (7,6,0), 73 => (0,0,14), 74 => (15,15,0), 75 => (6,6,0), 76 => (0,2,15), 77 => (0,1,15), 78 => (8,8,2), 79 => (6,6,0), 80 => (15,15,0), 81 => (2,1,2), 82 => (0,0,15), 83 => (15,15,0), 84 => (6,6,0), 85 => (0,1,15), 86 => (15,15,0), 87 => (6,6,0), 88 => (0,0,8), 89 => (0,0,15), 90 => (15,15,0), 91 => (10,10,0), 92 => (15,15,0), 93 => (2,2,3), 94 => (0,1,15), 95 => (1,3,14), 96 => (0,1,14), 97 => (0,1,14), 98 => (0,1,14), 99 => (1,3,14), 100 => (0,1,14), 101 => (0,1,14), 102 => (0,1,14), 103 => (1,3,14), 104 => (0,1,14), 105 => (1,3,14), 106 => (0,1,14), 107 => (0,1,14), 108 => (0,1,14), 109 => (0,1,14), 110 => (1,3,14), 111 => (0,1,14), 112 => (0,2,14), 113 => (0,1,14), 114 => (0,1,14), 115 => (1,3,14), 116 => (0,1,14), 117 => (0,1,14), 118 => (0,1,14), 119 => (1,3,14), 120 => (0,1,14), 121 => (0,1,14), 122 => (0,1,14), 123 => (1,3,14), 124 => (0,1,14), 125 => (0,1,14), 126 => (0,1,14), 127 => (1,3,14), 128 => (0,1,14), 129 => (0,1,14), 130 => (0,1,14), 131 => (1,3,14), 132 => (0,1,14), 133 => (0,1,14), 134 => (0,1,14), 135 => (1,3,14), 136 => (0,1,14), 137 => (0,1,14), 138 => (0,1,14), 139 => (1,3,14), 140 => (0,1,14), 141 => (0,1,14), 142 => (0,1,14), 143 => (1,3,14), 144 => (0,1,14), 145 => (0,1,14), 146 => (0,1,14), 147 => (1,3,14), 148 => (0,1,14), 149 => (0,1,14), 150 => (0,1,14), 151 => (1,3,14), 152 => (0,1,14), 153 => (0,1,14), 154 => (0,1,14), 155 => (1,3,14), 156 => (0,1,14), 157 => (0,1,14), 158 => (0,1,14), 159 => (1,3,14)), 
			99 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,1,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,1,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,1,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,1,14), 20 => (0,2,14), 21 => (0,1,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,1,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,1,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,1,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,1,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,1,14), 44 => (0,1,14), 45 => (0,1,14), 46 => (0,1,14), 47 => (1,3,14), 48 => (2,4,14), 49 => (1,3,14), 50 => (1,3,14), 51 => (0,2,14), 52 => (2,3,12), 53 => (8,0,0), 54 => (8,0,0), 55 => (4,4,12), 56 => (3,6,14), 57 => (7,8,14), 58 => (0,2,14), 59 => (2,4,14), 60 => (0,2,14), 61 => (4,6,14), 62 => (4,5,5), 63 => (7,6,0), 64 => (8,8,0), 65 => (0,0,5), 66 => (1,3,14), 67 => (4,6,14), 68 => (6,8,14), 69 => (1,3,15), 70 => (8,7,0), 71 => (2,2,0), 72 => (1,4,15), 73 => (0,3,15), 74 => (7,7,0), 75 => (7,7,0), 76 => (9,8,0), 77 => (3,3,0), 78 => (3,3,0), 79 => (0,0,15), 80 => (8,7,0), 81 => (3,3,0), 82 => (0,1,15), 83 => (8,7,0), 84 => (3,3,0), 85 => (0,1,15), 86 => (7,7,0), 87 => (7,7,0), 88 => (9,8,0), 89 => (3,3,0), 90 => (7,7,0), 91 => (2,2,3), 92 => (7,7,0), 93 => (3,3,0), 94 => (0,1,15), 95 => (0,1,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,1,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,1,14), 104 => (0,2,14), 105 => (0,1,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,1,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,1,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,1,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,1,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,1,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,1,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,1,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,1,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,1,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,1,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,1,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,1,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,1,14)), 
			100 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,1,14), 48 => (0,1,14), 49 => (0,1,14), 50 => (0,1,14), 51 => (1,3,14), 52 => (0,1,14), 53 => (0,4,15), 54 => (2,5,15), 55 => (0,2,14), 56 => (2,4,14), 57 => (0,1,14), 58 => (1,3,14), 59 => (5,8,14), 60 => (0,1,14), 61 => (6,8,14), 62 => (3,5,14), 63 => (0,2,15), 64 => (2,4,15), 65 => (1,3,14), 66 => (0,2,14), 67 => (1,3,14), 68 => (1,3,14), 69 => (0,1,14), 70 => (0,1,15), 71 => (0,1,15), 72 => (0,1,14), 73 => (0,1,14), 74 => (0,1,15), 75 => (0,1,15), 76 => (0,1,15), 77 => (0,1,15), 78 => (0,1,15), 79 => (0,2,14), 80 => (0,1,15), 81 => (0,1,15), 82 => (0,2,14), 83 => (0,1,15), 84 => (0,1,15), 85 => (0,2,14), 86 => (0,1,15), 87 => (0,1,15), 88 => (0,1,15), 89 => (0,1,15), 90 => (0,1,15), 91 => (0,1,15), 92 => (0,1,15), 93 => (0,1,15), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			101 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,1,14), 51 => (1,3,14), 52 => (1,3,14), 53 => (0,2,14), 54 => (0,1,14), 55 => (1,3,14), 56 => (2,4,14), 57 => (0,2,14), 58 => (1,3,14), 59 => (0,2,14), 60 => (1,3,14), 61 => (1,3,14), 62 => (2,4,14), 63 => (0,1,14), 64 => (0,2,14), 65 => (2,4,14), 66 => (0,1,14), 67 => (0,2,14), 68 => (1,3,14), 69 => (0,1,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			102 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,1,14), 52 => (0,1,14), 53 => (0,1,14), 54 => (0,2,14), 55 => (0,1,14), 56 => (0,1,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,1,14), 62 => (1,3,14), 63 => (1,3,14), 64 => (0,1,14), 65 => (0,1,14), 66 => (0,2,14), 67 => (0,1,14), 68 => (0,1,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			103 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,1,14), 58 => (0,1,14), 59 => (0,1,14), 60 => (0,2,14), 61 => (0,1,14), 62 => (0,1,14), 63 => (0,1,14), 64 => (0,1,14), 65 => (0,1,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,1,14), 71 => (0,1,14), 72 => (0,1,14), 73 => (0,2,14), 74 => (0,1,14), 75 => (0,1,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,1,14), 80 => (0,1,14), 81 => (0,2,14), 82 => (0,1,14), 83 => (0,1,14), 84 => (0,1,14), 85 => (0,1,14), 86 => (0,1,14), 87 => (0,1,14), 88 => (0,1,14), 89 => (0,1,14), 90 => (0,1,14), 91 => (0,1,14), 92 => (0,1,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,1,14), 99 => (0,1,14), 100 => (0,1,14), 101 => (0,1,14), 102 => (0,1,14), 103 => (0,1,14), 104 => (0,1,14), 105 => (0,1,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,1,14), 113 => (0,1,14), 114 => (0,1,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,1,14), 121 => (0,1,14), 122 => (0,1,14), 123 => (0,2,14), 124 => (0,1,14), 125 => (0,1,14), 126 => (0,1,14), 127 => (0,2,14), 128 => (0,1,14), 129 => (0,1,14), 130 => (0,1,14), 131 => (0,2,14), 132 => (0,1,14), 133 => (0,1,14), 134 => (0,1,14), 135 => (0,1,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,1,14), 141 => (0,1,14), 142 => (0,1,14), 143 => (0,1,14), 144 => (0,1,14), 145 => (0,1,14), 146 => (0,1,14), 147 => (0,1,14), 148 => (0,2,14), 149 => (0,1,14), 150 => (0,1,14), 151 => (0,1,14), 152 => (0,2,14), 153 => (0,1,14), 154 => (0,1,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			104 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,1,14), 61 => (0,1,14), 62 => (8,9,14), 63 => (7,8,14), 64 => (7,8,14), 65 => (2,3,12), 66 => (0,1,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,1,14), 70 => (7,8,14), 71 => (7,8,14), 72 => (7,8,14), 73 => (0,0,13), 74 => (8,9,14), 75 => (3,4,13), 76 => (0,1,14), 77 => (0,2,14), 78 => (0,0,14), 79 => (8,9,14), 80 => (1,2,11), 81 => (0,1,14), 82 => (8,9,14), 83 => (2,3,13), 84 => (7,8,14), 85 => (3,4,13), 86 => (7,8,14), 87 => (7,8,14), 88 => (8,9,14), 89 => (3,4,13), 90 => (7,8,14), 91 => (7,8,14), 92 => (7,8,14), 93 => (0,0,13), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,1,14), 98 => (8,9,14), 99 => (2,3,13), 100 => (7,8,14), 101 => (3,4,13), 102 => (2,4,14), 103 => (7,8,14), 104 => (8,9,14), 105 => (4,5,13), 106 => (0,1,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,1,14), 112 => (3,5,14), 113 => (8,7,12), 114 => (9,8,12), 115 => (0,0,13), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,1,14), 120 => (4,5,14), 121 => (7,8,14), 122 => (3,4,13), 123 => (0,1,14), 124 => (2,4,14), 125 => (8,9,14), 126 => (7,8,14), 127 => (0,0,13), 128 => (2,4,14), 129 => (8,9,14), 130 => (7,8,14), 131 => (0,0,13), 132 => (8,9,14), 133 => (7,8,14), 134 => (7,8,14), 135 => (2,3,12), 136 => (0,1,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,1,14), 140 => (3,4,14), 141 => (7,8,14), 142 => (8,9,14), 143 => (3,4,13), 144 => (7,8,14), 145 => (7,8,14), 146 => (8,9,14), 147 => (4,5,13), 148 => (0,0,14), 149 => (8,9,14), 150 => (8,9,14), 151 => (3,4,13), 152 => (0,0,14), 153 => (8,9,14), 154 => (1,2,11), 155 => (0,1,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			105 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,1,14), 62 => (5,5,11), 63 => (6,6,12), 64 => (15,15,14), 65 => (6,6,11), 66 => (0,1,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,0,14), 70 => (15,15,14), 71 => (4,4,12), 72 => (15,15,14), 73 => (7,6,12), 74 => (15,15,14), 75 => (7,7,12), 76 => (0,1,14), 77 => (0,1,14), 78 => (3,4,14), 79 => (12,12,13), 80 => (10,10,12), 81 => (0,0,13), 82 => (14,14,14), 83 => (5,5,12), 84 => (15,15,14), 85 => (1,1,12), 86 => (15,15,14), 87 => (11,11,13), 88 => (3,2,12), 89 => (0,0,12), 90 => (15,15,14), 91 => (4,4,12), 92 => (15,15,14), 93 => (8,7,12), 94 => (0,1,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,0,14), 98 => (15,15,14), 99 => (5,5,12), 100 => (15,15,14), 101 => (6,6,12), 102 => (13,12,13), 103 => (12,12,13), 104 => (6,6,12), 105 => (0,0,12), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,1,14), 112 => (8,7,12), 113 => (11,11,12), 114 => (1,1,12), 115 => (9,9,12), 116 => (0,1,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,0,14), 121 => (15,15,14), 122 => (7,7,12), 123 => (0,0,14), 124 => (15,15,14), 125 => (5,5,12), 126 => (15,15,14), 127 => (6,5,12), 128 => (15,15,14), 129 => (5,5,12), 130 => (15,15,14), 131 => (7,6,12), 132 => (4,4,11), 133 => (6,6,12), 134 => (15,15,14), 135 => (6,6,11), 136 => (0,1,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,0,14), 140 => (14,13,13), 141 => (12,12,13), 142 => (6,6,12), 143 => (0,0,12), 144 => (15,15,14), 145 => (11,11,13), 146 => (3,2,12), 147 => (0,0,12), 148 => (13,13,14), 149 => (6,6,12), 150 => (6,6,12), 151 => (2,2,12), 152 => (2,4,14), 153 => (12,12,13), 154 => (10,10,12), 155 => (0,0,13), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			106 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,0,14), 62 => (15,15,14), 63 => (7,6,12), 64 => (0,0,12), 65 => (0,0,13), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,0,14), 70 => (15,15,14), 71 => (11,11,13), 72 => (7,7,12), 73 => (0,0,13), 74 => (15,15,14), 75 => (7,6,12), 76 => (0,0,14), 77 => (0,1,14), 78 => (8,9,13), 79 => (6,6,12), 80 => (15,15,14), 81 => (1,1,11), 82 => (0,0,14), 83 => (15,15,14), 84 => (6,6,12), 85 => (0,0,14), 86 => (15,15,14), 87 => (6,6,12), 88 => (0,0,12), 89 => (0,0,14), 90 => (15,15,14), 91 => (10,10,13), 92 => (15,15,14), 93 => (2,2,12), 94 => (0,1,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,0,14), 98 => (13,13,14), 99 => (5,5,12), 100 => (15,15,14), 101 => (2,2,12), 102 => (0,0,13), 103 => (0,0,12), 104 => (15,15,14), 105 => (8,8,12), 106 => (0,1,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,1,14), 112 => (8,8,12), 113 => (5,5,11), 114 => (8,8,13), 115 => (3,3,12), 116 => (0,1,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,0,14), 121 => (15,15,14), 122 => (7,6,12), 123 => (0,1,14), 124 => (1,2,12), 125 => (6,6,12), 126 => (15,15,14), 127 => (7,7,12), 128 => (0,1,12), 129 => (6,6,12), 130 => (15,15,14), 131 => (6,5,12), 132 => (15,15,14), 133 => (7,6,12), 134 => (0,0,12), 135 => (0,0,13), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,0,13), 141 => (0,0,12), 142 => (15,15,14), 143 => (7,6,12), 144 => (15,15,14), 145 => (6,6,12), 146 => (0,0,12), 147 => (0,0,14), 148 => (15,15,14), 149 => (5,5,12), 150 => (15,15,14), 151 => (7,6,12), 152 => (7,8,13), 153 => (6,6,12), 154 => (15,15,14), 155 => (1,1,11), 156 => (0,1,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			107 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,1,14), 62 => (7,7,12), 63 => (7,7,12), 64 => (9,8,12), 65 => (4,3,12), 66 => (0,1,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,1,14), 70 => (8,7,12), 71 => (3,2,11), 72 => (0,1,14), 73 => (0,1,14), 74 => (7,7,12), 75 => (7,7,12), 76 => (9,8,12), 77 => (3,3,12), 78 => (3,3,12), 79 => (0,0,14), 80 => (8,7,12), 81 => (4,3,12), 82 => (0,1,14), 83 => (8,7,12), 84 => (3,3,12), 85 => (0,1,14), 86 => (7,7,12), 87 => (7,7,12), 88 => (9,8,12), 89 => (3,3,12), 90 => (7,7,12), 91 => (2,2,12), 92 => (7,7,12), 93 => (3,3,12), 94 => (0,1,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,0,14), 99 => (9,8,12), 100 => (2,2,12), 101 => (0,0,14), 102 => (9,8,12), 103 => (8,8,12), 104 => (7,7,12), 105 => (0,0,13), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,0,13), 113 => (9,8,12), 114 => (3,3,12), 115 => (0,1,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,1,14), 120 => (4,5,13), 121 => (7,7,12), 122 => (8,8,12), 123 => (0,0,12), 124 => (9,8,12), 125 => (7,7,12), 126 => (7,7,12), 127 => (0,0,13), 128 => (9,8,12), 129 => (7,7,12), 130 => (7,7,12), 131 => (0,0,13), 132 => (7,7,12), 133 => (7,7,12), 134 => (9,8,12), 135 => (4,3,12), 136 => (0,1,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,1,14), 140 => (9,8,12), 141 => (8,8,12), 142 => (7,7,12), 143 => (0,0,13), 144 => (7,7,12), 145 => (7,7,12), 146 => (9,8,12), 147 => (3,3,12), 148 => (2,2,12), 149 => (8,8,12), 150 => (7,7,12), 151 => (3,2,12), 152 => (3,3,12), 153 => (0,0,14), 154 => (8,7,12), 155 => (4,3,12), 156 => (0,1,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			108 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,1,14), 63 => (0,1,14), 64 => (0,1,14), 65 => (0,1,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,1,14), 71 => (0,1,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,1,14), 75 => (0,1,14), 76 => (0,1,14), 77 => (0,1,14), 78 => (0,1,14), 79 => (0,2,14), 80 => (0,1,14), 81 => (0,1,14), 82 => (0,2,14), 83 => (0,1,14), 84 => (0,1,14), 85 => (0,2,14), 86 => (0,1,14), 87 => (0,1,14), 88 => (0,1,14), 89 => (0,1,14), 90 => (0,1,14), 91 => (0,1,14), 92 => (0,1,14), 93 => (0,1,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,1,14), 100 => (0,1,14), 101 => (0,2,14), 102 => (0,1,14), 103 => (0,1,14), 104 => (0,1,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,1,14), 114 => (0,1,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,1,14), 121 => (0,1,14), 122 => (0,1,14), 123 => (0,2,14), 124 => (0,1,14), 125 => (0,1,14), 126 => (0,1,14), 127 => (0,2,14), 128 => (0,1,14), 129 => (0,1,14), 130 => (0,1,14), 131 => (0,2,14), 132 => (0,1,14), 133 => (0,1,14), 134 => (0,1,14), 135 => (0,1,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,1,14), 141 => (0,1,14), 142 => (0,1,14), 143 => (0,2,14), 144 => (0,1,14), 145 => (0,1,14), 146 => (0,1,14), 147 => (0,1,14), 148 => (0,1,14), 149 => (0,1,14), 150 => (0,1,14), 151 => (0,1,14), 152 => (0,1,14), 153 => (0,2,14), 154 => (0,1,14), 155 => (0,1,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			109 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			110 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)), 
			111 => (0 => (0,2,14), 1 => (0,2,14), 2 => (0,2,14), 3 => (0,2,14), 4 => (0,2,14), 5 => (0,2,14), 6 => (0,2,14), 7 => (0,2,14), 8 => (0,2,14), 9 => (0,2,14), 10 => (0,2,14), 11 => (0,2,14), 12 => (0,2,14), 13 => (0,2,14), 14 => (0,2,14), 15 => (0,2,14), 16 => (0,2,14), 17 => (0,2,14), 18 => (0,2,14), 19 => (0,2,14), 20 => (0,2,14), 21 => (0,2,14), 22 => (0,2,14), 23 => (0,2,14), 24 => (0,2,14), 25 => (0,2,14), 26 => (0,2,14), 27 => (0,2,14), 28 => (0,2,14), 29 => (0,2,14), 30 => (0,2,14), 31 => (0,2,14), 32 => (0,2,14), 33 => (0,2,14), 34 => (0,2,14), 35 => (0,2,14), 36 => (0,2,14), 37 => (0,2,14), 38 => (0,2,14), 39 => (0,2,14), 40 => (0,2,14), 41 => (0,2,14), 42 => (0,2,14), 43 => (0,2,14), 44 => (0,2,14), 45 => (0,2,14), 46 => (0,2,14), 47 => (0,2,14), 48 => (0,2,14), 49 => (0,2,14), 50 => (0,2,14), 51 => (0,2,14), 52 => (0,2,14), 53 => (0,2,14), 54 => (0,2,14), 55 => (0,2,14), 56 => (0,2,14), 57 => (0,2,14), 58 => (0,2,14), 59 => (0,2,14), 60 => (0,2,14), 61 => (0,2,14), 62 => (0,2,14), 63 => (0,2,14), 64 => (0,2,14), 65 => (0,2,14), 66 => (0,2,14), 67 => (0,2,14), 68 => (0,2,14), 69 => (0,2,14), 70 => (0,2,14), 71 => (0,2,14), 72 => (0,2,14), 73 => (0,2,14), 74 => (0,2,14), 75 => (0,2,14), 76 => (0,2,14), 77 => (0,2,14), 78 => (0,2,14), 79 => (0,2,14), 80 => (0,2,14), 81 => (0,2,14), 82 => (0,2,14), 83 => (0,2,14), 84 => (0,2,14), 85 => (0,2,14), 86 => (0,2,14), 87 => (0,2,14), 88 => (0,2,14), 89 => (0,2,14), 90 => (0,2,14), 91 => (0,2,14), 92 => (0,2,14), 93 => (0,2,14), 94 => (0,2,14), 95 => (0,2,14), 96 => (0,2,14), 97 => (0,2,14), 98 => (0,2,14), 99 => (0,2,14), 100 => (0,2,14), 101 => (0,2,14), 102 => (0,2,14), 103 => (0,2,14), 104 => (0,2,14), 105 => (0,2,14), 106 => (0,2,14), 107 => (0,2,14), 108 => (0,2,14), 109 => (0,2,14), 110 => (0,2,14), 111 => (0,2,14), 112 => (0,2,14), 113 => (0,2,14), 114 => (0,2,14), 115 => (0,2,14), 116 => (0,2,14), 117 => (0,2,14), 118 => (0,2,14), 119 => (0,2,14), 120 => (0,2,14), 121 => (0,2,14), 122 => (0,2,14), 123 => (0,2,14), 124 => (0,2,14), 125 => (0,2,14), 126 => (0,2,14), 127 => (0,2,14), 128 => (0,2,14), 129 => (0,2,14), 130 => (0,2,14), 131 => (0,2,14), 132 => (0,2,14), 133 => (0,2,14), 134 => (0,2,14), 135 => (0,2,14), 136 => (0,2,14), 137 => (0,2,14), 138 => (0,2,14), 139 => (0,2,14), 140 => (0,2,14), 141 => (0,2,14), 142 => (0,2,14), 143 => (0,2,14), 144 => (0,2,14), 145 => (0,2,14), 146 => (0,2,14), 147 => (0,2,14), 148 => (0,2,14), 149 => (0,2,14), 150 => (0,2,14), 151 => (0,2,14), 152 => (0,2,14), 153 => (0,2,14), 154 => (0,2,14), 155 => (0,2,14), 156 => (0,2,14), 157 => (0,2,14), 158 => (0,2,14), 159 => (0,2,14)) 

		)
	);
	
	BEGIN	
		
	-- Processo de controle do HSync
	PROCESS(CLOCK_27(0))
		BEGIN
		IF(CLOCK_27(0)'EVENT and CLOCK_27(0) = '1') THEN
			-- ========================================
			--   parte do controle externo das imagens
			-- ========================================
			showDisplay <= (enableHS and enableVS) ='1';
			showColor <= '1'; --(enableHS and enableVS);
			hideColor <= '0';
			
			-- ========================================
			--   parte do controle do desenho
			-- ========================================
			quadrado <= (xInit <= drawHS and drawHS < xEnd and yInit <= drawVS and drawVS < yEnd);
					
			-- constrole de contagem
			IF (countHS < 809) THEN
				countHS <= countHS + 1;
			ELSE
				countHS <= 0;
			END IF;
			
			-- controle do Sincronismo
			IF (0 <= countHS and countHS <= 102) THEN
				VGA_HS <= '0';
			ELSE
				VGA_HS <= '1';
			END IF;
		
			-- controle do enable do HSync : 640 px (793 - 153 = 640)
			IF ( 153 <= countHS and countHS < 793 ) THEN
				enableHS <= '1';
			ELSE
				-- testar consistencia do startdraw
				-- drawHS <= 0;
				enableHS <= '0';
			END IF;

		END IF;
	END PROCESS;

	
	
	-- Processo de controle do hSinc
	PROCESS (VGA_HS)
		BEGIN
		IF (VGA_HS'EVENT and  VGA_HS = '1') THEN
			-- constrole de contagem
			IF (countVS < 525) THEN
				countVS <= countVS + 1;
			ELSE
				countVS <= 0;
			END IF;
			
			-- controle do Sincronismo
			IF (0 <= countVS and countVS <= 2) THEN
				VGA_VS <= '0';
			ELSE
				VGA_VS <= '1';
			END IF;
		
			-- controle do enable do HSync : 480 px (515-35 = 480)
			IF ( 35 <= countVS and countVS < 515 ) THEN
			
				enableVS <= '1';
			ELSE
				-- testar consistencia do start draw
				-- drawVS <= 0;
				enableVS <= '0';
			END IF;	
		
		END IF;
			
	END PROCESS;
	
	-- processo de desenhar o quadrado
	PROCESS (CLOCK_27(0))
	-- PROCESS (CLOCK_50)
		BEGIN
		-- obs
		-- showColor corresponte a operacao AND enableVS e enableHS avaliando bits quando estiverem ativos
		-- showDisplay corresponde operacao AND enableVS e enableHS em boleano
		IF (CLOCK_27(0)'EVENT and CLOCK_27(0) = '0') THEN

			IF(enableHS = '0') THEN
				drawHS <= 0;
				
			END IF;
			
			IF(enableVS = '0') THEN
				drawVS <= 0;
			END IF;
			
			
			IF (showDisplay) THEN
				IF (drawHS < 639) THEN
					drawHS <= drawHS + 1;
				ELSE
					IF (drawVS < 480) THEN
						drawVS <= drawVS + 1;
					ELSE
						-- drawVS <= 0;
					END IF;
					-- drawHS <= 0;
				END IF;


				-- IF (xInit <= drawHS and drawHS < xEnd ) and  (yInit <= drawVS and drawVS < yEnd) then
					-- VGA_R <= 15;
					-- VGA_G <= 0;
					-- VGA_B <= 15;
				-- else
					-- VGA_R <= 0;
					-- VGA_G <= 0;
					-- VGA_B <= 0;
				-- end if;
				IF not (
					(( 0 <= drawHS and drawHS < 159 ) and (0 <= drawVS and drawVS < 111)) or
					((xInit <= drawHS and drawHS < xEnd ) and  (yInit <= drawVS and drawVS < yEnd))
				) THEN
					VGA_R <= 0;
					VGA_G <= 0;
					VGA_B <= 15;
				END IF;
				
				IF ( 0 <= drawHS and drawHS < 159 ) and (0 <= drawVS and drawVS < 111) THEN
					VGA_R <= sonic(0)(drawVS, drawHS).r;
					VGA_G <= sonic(0)(drawVS, drawHS).g;
					VGA_B <= sonic(0)(drawVS, drawHS).b;
				END IF;
				
				
				IF (xInit <= drawHS and drawHS < xEnd ) and  (yInit <= drawVS and drawVS < yEnd) then
				-- IF (315 <= drawHS and drawHS < 325 ) and  (315 <= drawVS and drawVS < 325) then
					VGA_R <= pacman(pacmanFrame)(drawVS - yInit, drawHS - xInit).r;
					VGA_G <= pacman(pacmanFrame)(drawVS - yInit, drawHS - xInit).g;
					VGA_B <= pacman(pacmanFrame)(drawVS - yInit, drawHS - xInit).b;
				END if;
			ELSE
			
				
			-- eh obrigatorio manter o nivel logico em 0 quando nao for autorizado o desenho
			-- caso constrario nao eh projetado no display
				VGA_R <= 0;
				VGA_G <= 0;
				VGA_B <= 0;
				
				 
			END IF;
	
		END IF;
	
	END PROCESS;
	
	-- controle do processo de movimento
	PROCESS (CLOCK_27(0))
		BEGIN
		IF(CLOCK_27(0)'EVENT and CLOCK_27(0) = '0') THEN
			IF (not startController = '1') THEN
				startController <= '1';
				
				xInit <= 315;
				xEnd <= 325;
				
				yInit <= 235;
				yEnd <= 245;
				
				moveDelay <= 0;
				
				pacmanFrame <=0 ;
			ELSE
				IF ((KEY(3) OR KEY(2) OR KEY(1) OR KEY(0)) = '1' )THEN 
					IF (moveDelay < tempo) THEN
						moveDelay <= moveDelay + 1;
						
					ELSE
						moveDelay <= 0;
					END IF;

					
				END IF;
				
				-- cima
				IF (KEY(3) = '0') THEN
					IF (yInit > 0 and moveDelay = tempo) THEN
						yInit <= yInit - 1;
						yEnd <= yEnd - 1;
											
						IF (pacmanFrame < 4) THEN
							pacmanFrame <= pacmanFrame + 1;
						ELSE
							pacmanFrame <= pacmanFrame + 0;
						END IF;
						
					END IF;
					
					LEDG(5) <= '1';
				ELSE
					LEDG(5) <= '0';
				END IF;	
			
				-- baixo
				IF(KEY(2) = '0') THEN
					IF (yEnd < 480 and moveDelay = tempo) THEN
						yInit <= yInit + 1;
						yEnd <= yEnd + 1;
											
						IF (pacmanFrame < 4) THEN
							pacmanFrame <= pacmanFrame + 1;
						ELSE
							pacmanFrame <= pacmanFrame + 0;
						END IF;
						
					END IF;
					LEDG(7) <= '1';
				ELSE
					LEDG(7) <= '0';
				END IF;

				
				-- esquerda
				IF (KEY(1) = '0') THEN
					IF (xInit > 0 and moveDelay = tempo) THEN
						xInit <= xInit - 1;
						xEnd <= xEnd - 1;
											
						IF (pacmanFrame < 4) THEN
							pacmanFrame <= pacmanFrame + 1;
						ELSE
							pacmanFrame <= pacmanFrame + 0;
						END IF;
						
					END IF;
					LEDG(3) <= '1';
				ELSE
					LEDG(3) <= '0';
				END IF;	
				
				-- direita
				IF (KEY(0) = '0') THEN
					IF (xEnd < 640 and moveDelay = tempo) then
						xInit <= xInit + 1;
						xEnd <= xEnd + 1;
											
						IF (pacmanFrame < 4) THEN
							pacmanFrame <= pacmanFrame + 1;
						ELSE
							pacmanFrame <= pacmanFrame + 0;
						END IF;

					END IF;
					LEDG(1) <= '1';
				ELSE
					LEDG(1) <= '0';
				END IF;
				
			END IF;
		
		END IF;
	
	END PROCESS;
	
END Kim;